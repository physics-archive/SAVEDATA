MPQ    �Z	    h�  h                                                                                 �L=|�����d@�|K��}�C�P`�}�h�"ä�,��H!bogm�L�!0�<5��!6�X���q�֬��U����.%C�90Ì�/�3z������4D�g��E9���i��"�^�glnl4��4 x�@��l5�0dZ��vx�8��O���Gm�n	#q�K��G#R�ѿk9A4nd��*c�8Yo�7�����4�Ǆ0$�&��ҏ����H��e92��ZZ�E��{�E��&c�C��o��w��c�C�{kl�Yt�Q���s��F�Ө�r�1���
2�	|�i����h�?x� 1g6�!��=��/ߠ��2�s�nG�|�;�Gs�${�MmY��\�	A�Sk�1Qx�)�dK[z���L��	��o�)��_��A)�I�8�QPpOy?AF����S���
�j�F��9�#�\<@xKc����y��C�l��>�+�"'	6%��%t#քr��(���[��Z�P�*7۷f�,�ݞ(C�qo�u�s����/i�O+di���S���fD #�*C��3"���=����i+B�"D�#"t�Xr�_f��vU��=WZh��1��o� �(綠M���
3�g@_��L�����"Ùl�vY]4Sp��l��]�"��m豳i0��K��E�ub'����/��r� ����L\�բ� ����<p%Մ�yl?�Hu�g�ΪmW}�+*��P���]5a�HoggDuxK�䏟�8�K���v��~3�:�J�i��<��[�:A�Lq4Ȧh��t�(	����8u:n�C��j�g�W�@U{6s������f� �FdF����i=�a�9t�#uV)��qv�AZM��;�~�\��y�ܷ�z�����wv�R�޴3M^�����B�<~��-cU�Kb�ǃP����g�^�5�Z��c�XIA&�9���[���.'�)8�.F����}o�oQ����`�DrO�蟭�&%��6ǈ"��|�V�0��R�#�U�[�e-���S��
��Y��;Z�Q;UCV<3_�@-/��'
�	.4��CG�P�){��ǋ8�'�'*,�]���W��7���k�.��1�U��3������n��`0A<EL�W�^���kHe�:S㚳�D���g@����T�����6���b])Z/���Tw��mʤJ�[�[����r�er:Rmm4��N|oN�%%��|u<��~��/�PD�r��c��*�?�16�3�6�lr�l��k��	���QB5R=�=AO���>���/>ߍ����V��7��E��X���T�|@�5���a��s̻��Ԏn�;J]��y�o��}ݱ���D���9U�sd��������'t��z�<޶��ej�!�P�ۻC�wO�0BG�,�R���fy�]�qRs̓Z��f��:">��Q���(K�ϓ�~��7�b�7\�����P]�&��B��R����=�U[�#���� �~��G��h^s�Q��I*Yk-��>�u{�&Q�)�~���)�ap�f{=pb�_w�J��:$59���'*<�fޝ�rb�3N\�k�?�͠�'�?���VK?)`Ι!
�C!F�J��Ϳ�x���?�W��9���̞�.H���7���E�@�ȏ�����(>ӱ1��L�@uC��W�Aȸ]Ɵ�1��#/dk��a������5Տ����쉚w!su/�0^U����n2 �mw�0Jm���<���hSڷ���g>řj��ki���}��!t��p��H���������Ո�{���_˱JO�6/ggP� �|&	��Q�8|sE�l�|�<_�aS������W �9[�n�󂈍U�D�h���d�!I�jaR�^:(���i�Ȇ��h�Z���,Q�'W"���Ƶ��N�Tv.��] ���4P|=��_'7�
��Sl��hu�^P����ˀ�-Tq�@���<`���iy��G0�ٙs�À`v�E2+	�aX7����g�b盙s�,�v���s����0����m|@1���b-}��E�M��kTk���/��.�W�]n��BRa0G$Y��{�RN}�h
D#~9��'׬ѣ��`Xq8*�.zx��~oBM@�)��E ����?:ovt�%I�&C��{�n�������w��`[ �b9��<1�>S�Ȳ&����d��� ��cŕg~ˈI�ܕ�mXnG �䥢(
�����6���N8<���l���S�jɵ�kp�l�R�"[�3B�w"|�		Z�+�F��P,����c�ć"A�?�!�M�C0�u��9}#��7<���n`��UC&e6���1�1�+Ȼ���ୠ`�>��i�����%�(p� $��I}����Wf�_��-��#����}��L�]����U��ۨ�op���z����:��V�O�����eh�Ax\YSt���ݱO�3�ϹP��!��D�,j�������7�0��c�1ћy�d����Ƙ�i�)-=�ꥇt{G6�c����� ��xD��"����=Q�P`��L��ڻ7���:P��푳LII��{GB8.q(���$�����n�<�H�I|��GcւN};7Ye��r��A]XmP{���Q�B��(ld�$����qe^Hi������^X����Ik�8�m`۟�ǁ�}m4&���s-���v uU��S��S>J�݆h�5@iRS�<)��2��:0k �@���sek��I
��A�v�c�76�A��Ѣk!�ſTl�w�PYz{��hg��WՆ�$�-�����C"��^��=0��+ˁ c�K�;['؛���3b�Cu��!���@\�;����A�*�k�J{ʗC��O[�O1���L"�@��/xl��%��9d�!e�=��6np�':c�*T;#��D	������x���k�{��.H
��1\�����ƿ�o:d�'-E		�����p���XTe��_�ZȑpD�gv�fϽ'?�۸�Ry �uU�D��N��yOV�pG�(�7��_n����$
z��E�Jk�G9�^��hᠭ�t�j��O���5o=J�ߵ6F
WǸ̪��8��PK�/w���s��yMn`W`w\(~��Kө�vơG����"?����Re ��@|R��]ܹ���L\����۷"7��K/&Z0�ӧ�`�m?z���ms�<�%�38[��4ߜ���A&��xy�O��X��nS%*��YjW��N����S��y�$�A���p�8�n����eo"���Zv���[�EW�4cٖZ�������Z����C6{&��Y�p�Q��s�F�9_Sb1ȑ�etT��Zi_B��Icx���gV�ż�c=�I��4�2_�nb�
wAE;�ws ����#���&�d
�S�_91l�)��	K6
��Y��繙	�������_�
.ADiԳ�_PK�R?|+���F�s	�r��
�u�F�N ��5��_K����!q��>�{�3��+r��	Qr��#�����#�x��U�`��7����r���(M���su��|���R����
׋�����T��A��#$<��bl���
X{$b��=R�ٞ�%�3^Κ������	$!W�P������*�k�� �<����Mw,���gxa��l�y� ꣥7�t�V���i]��p�kl�d���ʹ2<��.UӾMr���b����@�/A�� ��ȕ\S�#��`���&%pԀ���?���T����}Ft"�����G�5��FHju�D�E����/ȓ��'G�Q̥~n_4:[p�i���P�d��D7�g��4C����P��cr��pju57��jH�Ȧr��U��6s�ᔫ�ykUbT ޵���c�i5�i4��af�W��&�Vd�ݙAU��ߖ��*sy�R;:j����w�D��y�tMY�?�<F�B�m~'-�_�K=$��H��B�Y�W���Gc;AA&�9H*[���.b�`���m)���toAHEQ)�g�:�<`���O�H����%�+���GDM�V�56>�#���[9��O\��;�̴�;::V(���3:�uh���*�<�Gs7�)��˼B8��s'e�Ӆ��������������.��fݕ���u�3�,���7�i�����Az�r,L�u�N�u5�N����Jg��3���1��R[Q��s��	�]�� �� ywI��_]�v,���V�M��2m4�����|ʠ;��ɗʶ�5w��	���G�r\����?�����ه��ljs�Լ��8`(5���8ʺO����f�Ji^�m������r��E���X��aT�O���T��Ě���L��j�L����J��AyȎ[qW�8�s��hD��[���ɯ�������Y'Ϯ	z���'�e��?�+^Ȼ@}�W0=�&, ���̏�y�4q�-��5��f��"�RQă������p��{
��.��,<��Vm�]�q���X�REu-�A�=ek [����R���@��]C'>�s�SQ61>I��>k��>��5��~�)�_��f��a.����aXp=�[_�񸽗�`54���tR�*��"f�o�53)�qk����;�����F�U�K�`�){'!�p�C�,�3�FҲ;Ժ���%WF89�����Hp��7@Ll���թ�S4^���>��)�|K��5C�R$��Y(�X����#�&jȯ8�l���"�p}W��N>��,�w|u/�~�p �Y� �%>���m1
n��i�:��rf �W�^t�F̉Ȯ�}�3-�����s���H�b��\�W��ƶuق�O��N�O�!"V���w|��E��	��sP�E�
�w�D_)U�<���G��/���<�gU6�h�z�d�T�%fٱy֏�T��ˣ�ޞS�Z��G�'�''�&�ߛV����KT��8��*������7 :���:����u\���Ke˻I-�x�@��i<a���O�ޤ��T�����xvZ�_2�{LaS���XSj��K,I��.ɗ���S��mw����b�8q�y�M�ck/�a��P����1�I_���-aKehY\h�{�N��
�։9�����j��2 qS3���[���o}���Ŀ:E��%��:���v.h�%�v@C���{ϰ2�xv�{N&�A�[�l�9���1l|S��u&9���È9��L�g9>�I �9��DXI��G;5��=����п4�g��5NS����$��`�S���I6��g��}8�3�Ps=g	���+�Y����>�(	���}I�?���!���� 0�3�}���2�K����v&��L�KE��_�9+@��"��[y����aG���B����4���y�Y��R�_Df4u����B����'���Ε�UG��ֽ{oj$m����1��q@�*@�)�e0�xW9�tc�!�|7�N����~��̮�!j�?J��:w7;���)Ѷ��dxf�XϤu|-�Ք���iG�� �����b��?����[�V�=��P[��L�9���?��ȑ�3�'_F�M�B��q4��_�жE��<v< ��$=e����q�}6���r��Ю6��]�I@{�/ӳ��s��](g�$i�B�T̆q��i3�d�Z�s^���(RIf4|��l���_T���Y��n���8h�7�ŲU��E���wJ��=��m�5�&FS�����:d��?e {C����!k��AI%�Asc��6)U��l]!��忯�)wL��Y�^��':/hB�WV󦵺	-��*�5��"�L�^�
��n�+��>c>W�֫�ؖ/�ԎE C0 �!ұ7�Eh;ب����ň��E�;���:O��1��[��V�@�R�/L��kL��3&�|Of��G65j�墹7���;^&�ߝD��b��-�P��Q����
��#$��l��&0��Oo��H'迡	�hS�o���w=Jp�e$%��U#��9f�"|�#I���Rۓ?0��ru�=��tȄ�4��+�y�C�>�bJ�u#��~z�!I�E\RG��'���S�@Mta��*��O��=�+(�1hW"��T���Ϝ�����y��M	t `�\��z˵}���ա�:���>͖�!JR ���g��ףM��jL�~���|ɷ]!���+�h�/����c�{�m��ދ��;�w-�%*��8V��4:���G���H#y*�ƛ3n���*y��Ye
������B���$�w9���_�sI6�~#�e���8_Z�^��[~E��.c�	���p�R���Ղ���{�3OY�[�Q�*�s�)FTf^�S"1�Q���Y2i*5��^�x[rg�ƹ�WD|=�(?�V�2g1n}mU�%�;Ϗvs[�Ճ�X��SM���S�t�1���)K)�"T�ڂ�	�tx�ߴ_y�aA_��.Z�P&�<?�0��8������
l�F
�n��-�	wK١����`�9�F���+-nV	l߭�&�#�����>̲AK�Pl��/7{<^�w��tc(����u!�~��%��L�P�Ţ7�#�I�k�u#_mQ������m�eC�߸��X�����4��վ���Ĺ[AW5g������C,��ȉ ���,�M[o� �gӢ��'��;����U�O:���ݸ]FGNp�8�lD{jۘ잹M+���әo=��k�bMő��J/l�/疃]�-��\��Pض-f�X�%D���?b�ؒ�b����&}��曊 Lӂ�
5���He�_D+3K�Z���Jx�A۽�,��~��%:���i�}����h㡂*�4��䰡l������u0���G�jPΦ�s�U	�bs�ZJ� ��}K �D���$ouiO��a�B���J�V����c�AP�E�񶋗��<y�tT����s�w����x-MT��
kB}f�~BY�-Y�UK�������Pb��T����c��A\X�9��[j7.�p��_��$�N�@̫o��_QD��J�`��gOB_E�%�z%���>��=JV� ��I�#k+e[t�D���\�،��K�;е�q9�$3�:��n� >��E揗�8G.>�)��*���U8��'��<�>$c����g��n.�b���4���V3*�o�*�٨dc���^�����K�u�ް7ߚ�P���vLg��dh7?&П���n��A�^]_����h9w�2������$�x���(l<�Jm�S����|%�뛀ɲ?����[�1G��jr��F���?]L���1O٢�l�of诏+�s��5�^�3sYOc���:�e���I���24���E$`
X�m+T<C�Í�}��н�xF��E�t����J�ry����1����α'!D����������х�I'*��zV/�B�e`�ʃݤ�{�z�rO08�,[d����y,�qH(���f
h�"t��Q�#
�BGاE���]-���假g�����]��9��"�R ���'�=�۷[�=�Q��=#����3Ns���QQ�I mk㼗>8bd�\��)�`���$��aI���\hp�c_킻�2��5/l��ϝH*�`1f�Th��3>�k/X���	���M�ܰ#�K���)���! C�Xbny��M���ǟHb4W�9�P�̔vTHKl�7{��{y6�@�� �l�>	0���9��$C�w� �S��烷#�	�������(Y�ES�F�����wח/k��%H���! ��T��m�D���7���=�-_�h�ŏq��!O���} �K���&���yv�7]���]�����^H�G`K��q�On]��dz�7�@|<+����D�E%���r��_�������
ڵ�/$V��U���fiU��h�4�dm�@���D���_��>��~č�?]ZP(~�";('K��V��|7Tl#���w�T?S��D���7{�ϊ����Eu��͓_���5�-���@���<�4�
���!�Ϻo�y��v���2a�aN�f���̷�h���/�,�-h�f	e�?�����mr��z|:b�_�,�8M�Z7k
W����qK}�/�E߃<�af��Y�i�{|P�N�h�
z��9�h�b��b$lqn\j$��z�o����_��E�#t�Or:�H�vI|�%?�C��{
|� x�v+Q�q�m[vt
9ۮ�1��rS�I&Y�?⚔+�0���rg��I;��܋�X$��Gv����y�\Կ���o��Nn�����x�2S Qʵ� ��bF'��53���Xܻ	��q+��#��(j��d��X��q�?�k!�E���0�$<L�}Y~�-Ĉ����`�N&�B�ƞ��:#G+>�e����V��GFn���(��{�hh�<�J�����M�_�0]����s��gq�	P�U��v���o��(�Z�ψ��������dd�e��&xR9�t����SgC�i�9�F���8���\Jj-���7ne?��lf�ѳ�d�69�|8W��P#-s�}�4G�;>�\���1*�n[U��t�ۑi=�G�PVAL=����� H�v����ӆ@>Bn)zq�_�E�ǋ�5��*i<{�c��̧��4j[}1W�rfC]�Q��]NF|{����ǋ�x�+(b�v$��F��
q���i��5�^�Ķ���Ia�;�#�=�E+���+Ґ�����ݬ��U���Q��Jx5� 56�S�60�cq�po vf��RXkyk�I@�%A�cpQ�6d�^��&!���
��w�Y�Ή좭�h��W�1;�U+-�S�ϐu+"�0o^�eL&-�+�}cK���qbؑ�z��H�C�n�!��6O;��j!��`d�@���̑O��1�+8�B�@�6_/�+��}MD�רG���6P�B�Yxt(;���zO���G׬�a�e�����%��]`�&A��]Ѽ��o�/'�Z^	�Z����[\R���e��j�P��&��ݡ�� �� ��n�]�Ru���ặ�/:���R�^Q-����P^ƾU1gz*D�@m�G��p�|8����t�w����ߊWt=��,��W}O��HV�!m�%ɳq
v�L�qM��!`�+\�j��p�i�#i-�=�ëz+��oR�b��ي��o�^����ZLRv�ȸc����xI��9/���IW���cm5߮�|qò��%���8Q��4��գl��vy�J��Kfnɵ*��Y`���5��H/���/$P��su���,R�n!e���C�4Z�g��| EMc��?� �m��7��>tT4�{��>Y�f�Q�syg�F�_�t�1�.��y�:x�iE+��ٜ.x6[�g��	����=�'�߱�?2�n�N�m*�;�#Fs��D��\������S>�1�|�)�j�K�g]n��]	�	��:�!_4j�Az\@ԩ� P�6?�U�ӿ����(=
'�pF%s����͞�K�̭W���4�ͼ�}+�CT	�lfWn#g��2z䲮�j�Kb�aW�76�G�ﴬ��'(� f�u��x���͏�p‎g��P���E����#�����=�����N{�/��sΙٔ���tF��G�$����W���@����|��a%� ����U��M��Z��8�g.�����V��e�*���'P�]�  p�%�l�q�Sw�h:�$�B�t����b�*x���b/�S>�Q&C�H�!\I.*ؑgǓu/%�ӧ���?���L����:}<ew�e��ӽ�52�<H`�D�@[�Z��eH=��� �2�~�{�:��i���k����49�4�|��٤����u+��T��j�x��sU�W�s��[����z ��u�|����ij��a\�����V�k"B
gAK[-�Lpb����y��1r�ob�w'�կ�^MOj���&B8��~]�-��hK������޾�O�o�k�_c��6Aw��9S�[E_�.�P�����wJ��#o�3�Q_V��0+�`j�ZO}J���E�%{WLǙ�P�NDVI�,uS#F�K[����T�U�����j��;�Q��.�Y�3�;���l»A����i��l#G�d�)̭��8p�8m�A'��Y�ٷ!����HNn�C .�K�݋Ж����3e���ųӨ_5�q�m���_�k������Y˚��-���gQ;�#��A��H�x��@D�]�w���Еw��������`��~��	�#�+m>����|��4�V^�����+ȸ�]yK���rU�|����?�	��d��ٽ��l`�E节�׮�P5#��.<�O�m��o.xހu�c��n�J��7�E��?X�T�V(�H2��&���_� 
M�W�J.^%y�,�'pϮ��BP!D�a ���#�$RTB�z�'�a�z�-�] �e�4���{q��Q�H4�03�z,��ʛB�y/CEq�(���fE�"��Q��(�ϧ 4��_��b˘��.��<��|`]�g��SqR��g�B�V=[l[\���h���%H��!�HVsDmQl�I�H�k�>s��9�)����e�Zb�adY��׎�p��_(4R��d"5*X��*	N*m7�f/Hb�V�3��$kj��qM������MKN�)�9�!{�uC����@���x�ʞ埣##W���9�y�~�H&c�7�С��e�OR�	�'��>$���r��j��CP���C��N���B�{#`��C��b|u���-��������w2�*/&z��jI�O�K a��L�mg����嬇�P���w!�H�
�@����>��}��b�������y(�Rx��Rܞ�f��,hK�␯����O� ����R�1|�=������XUE�!��m�_�̘��q��%�l��8뻗���3��Ul��h��d�ӛϓ��n��J���Y-�z��Z�,��'h����V�D�T��������t!�,��O�7�� ���2ЯuRߎ�:u��1v�-%��@��w<�m�ź��-�J��T�v�#�2���aI����������ķv,?�"�Aq�=�v����mmSj�l.b^ўG?�M1k����7��9��.n`���v�a�iYR��{W��N.�W
�I9}ib׽D9�6�q����_��v�o�R���\E�Uw����:@�(vd�<%�ŷC�(:{E��ݮ�e�q(���Y�[1�d9�́1b��Sb^,&�3��5�*��h�t�g���IV�m�Y�X���G�E�s���ꌋ*3�N���y5�S��S[�ȵ+a�]�[�3S�3ss��	z�J+u���	�^�;��.��3��?IZ]!+O��v=�0j�w�}�_�(�w�i����&���Ax��+y�؍Xcg�Q�(���:��|��d��]�����wWi��H��_����QW�;�����e��D*5U}d��G"o ����W���A�g��s��I:e9)�xMYwt�Y�rs��_k���۲����L�j�����n7ɯ����� Adn'6�W8��L-{q�x6�GG�����'iڅ���)��o�="�PQ¦L�/v�h+!�DБ� �����{O�B	bDq�������Fʩ�8�<�\����,�6},2vM�r!��l�e]�b{�g����Q(]�^$+��Esq��ei)[U�lz^	��R�2I\nw�~�� ���z=����e����o�Gn�U����YJJ3�j����5�2Sq���@����� q�����Zk4Y�I[+Ai��cK��6���r�!�ϻ�et�w�Z�Y�^m�A�h���W̏C��4?-�,`��m�"M4�^����+\+lc��+��#،Wn�Dl0C��"!^�x�;�:�=����_��;hҗT�O��1�|\Ľ�@�:�/H����x���2"	�nq6k�G�%O�Q;�ǝ!$��L}�� ������� ��ٷ��⻳�\["ѷ�RoKr6'^?	�l��e�6a���heZT�K9��jҘ��������I�*u&���� ���_��Y��y9�X���+������z��7�;�GJ:�7�����t�0���=���=��'�wW����.[�<+������L��~�M?�Z`l�\9t�+A۩>͡���Æ�Y�F�iR6ܖ��kWQ����ڹ#�L͍�ȓju����+��
/7�Â�����m�A�W#�����%`��8L��4�)��E��qy ����n�N*��Y[�r�_�V��a�3$�H��N}-��/��ؑe�H�jZF���.��E�J�cjOZ�[����+��a�ܑ{W{�Y���Q�'8sTŶF�xd0��1�c&�v�|���Hi`A��Tv�xd�g�ō{U=�F?�С2�ڰn�O��N;���s�!�չ�����u&�S��P1�h�)ځK��6���ڸ�p	��q��=3_�I�A�3��$��Pܶ@?-�<�n�Y�ɷ��u
�UF@5D���S6KO";���/�D(,+�9�	����#BD�m�P�I�b�Fx��,�7��҇�����(��[��uWk����q8�;����?�+��[*#�/��3�/�����z�U�?�<��(D���B�K�r�⣼��(6W����]�֐�ܡ� � ���MH���z�g�����?��qV)�w-9����b�3]|�)p�2:l��w�<S��iD����O�1�[b�oÑ�h/"+m��L�c�c\ċ��l'����%A�O�
Ez?�<�ޣ��}�ԛ@p����5ͼ{H[_�D�m˳�2��8n�7�o���~:e:,�iz�\aj��&ȡ��C4����W��n�A�#u&���.�jyƦ��~U��?s��ū���&� ����?)��B6i�A�a��ʃ}�VK1��QAF�pߧI�H�|y���8��Jq�wb�I�J�MJ~9�M��B�e~xG�-O?K�ԙ�<��{a�J�e���clyA�#9�[ �[.Q�ꕖ�r��`�or�`Qz���+�`EĝO�U;�[�/%va��w�u�V5���� #!��[��,��F�Ύ��ŋu;F�a/�=3ˡu���V������MH�G���)��`��QO8H�0'+�tk��3`��T����.�T���D�{In3��q�`�%�Z'���5Q(�\�è���u~#��&���D����g������\n��BNS��{��]�l���X�wZ!�ʐU�*��n�8����^ۆm��ۀ�V/|�W�\!����� ��8៶<qr�[����?��#���2vlۖ�e�;��J�5�S��)%�Ovi�*Bmޛ�����I���#�]EZ��X��T�`��V����n�H��rՎZ�XJ�iky�������i�б]�iD��t����_��l�u0>'��}z�O�xleV$��:.���/��0.�^,d1���ByJz*q>���p�f���"�>Q������姻�܉��#ț������n�'4�]����3Rvk�]�=�K[7c8��#�sH��_[8~�s�MsQ��fIDxk�r�>������)��wŮ��a<u�R��p΢#_c}�h]�5%d�ׅ��*(.;fJ�^�3��k����,��ۗ�fp�K	��)���!��0Ct��'v҃G2�@`���Ww�l9y�̊�*Hzv7��*������d�q�.�>?.C����E��C�����ٸI�봝�_#/?������W�U�!6�|����Mw�<�/�'�����A <s���m{����Kިڣ��<��Ņ���״1y��}V�q�w��<Q�4�]�m����zT�A�]�g��}�+���O$�S�4�m�J|�z�~���$��E[ݮ�h��_:�ڲmK�@�k�%m̻r���nŕU�h��d#G��V4Ǳ�j7��_�4�����!Z�+S���'�����Ŕ�"+�Tb�a��ǋ����������|71���?���M��u����:�l��-�O�@�P<r�:���p�/|��[��/��v��2��oaDG�i���NjA��_�,�dɨ�xv�$&�mhD 0}�b,ǞbңM}'k���rtd��l���ɛ����a�%Y��{2�Nia�
���9x���@��g�q��̀w��o.�͕ۀE����6R%:���v0%5�Cs�R{�7��I���lE�'{[���9�1�S=�&���������Ϣ�gjVIqσ܁��Xڹ"G��^�g����E�}�N������.XS���V�X"lĎ��3.����	��+PR~�<���o���w܇�"�?��!F:Ǵ�0E-���V}�`��#̂�\�U�֐�&��3ռ����r+������j�L������x��&L�Bk0�ֲFh�*@h�CNU_U�f��"���i����E�$�U`��Ǽ/o{���9���T����˻=��N�e��kxH��tt�%�ɜ����D�<oۍ�0]8jc&;����7$��O���n�d�7��2X��Ugm-����s^G�F���#��B�r�d򯣎�7��o=��PLc1L��T�#�י4�`�lǫ��`����?B��&q������[��f�<qN���?��3?�B�H}'S��c�r��®��]D��{i3v�=�v���(X��$zZ��qѮ?i��o����^DIw�WIW;/��Q������i��=�@��D*��r�U�(����J�7�ԛ5,*SL���{(�.� l����k�f�Iv��A�Xcc&!H6�N!�=MB!��p��aw}�Y�9��/hӪ%W���zK-�%��F�"XY^)|{
�+7�Zc�y�ŧ]�؇~ԟ�8Ca�3!#�2,��;i�{x)�ʖ{��6������OG�1����8��@n^)/�4:�<�
sᔧ����)6�6����=*��;ŕ��Ȱ�q��>ʄ���!��{�.�1�q:���Ѳ�[o�a]'�C	��;������P�e�V�F�S�(L�SM��g��/�$O�e�u��8�צ*��v�\J0єA����e�4��˽�z`�#�6�{G�����.��it�v�-� ��=�咵"�)W3f⪅5�W	��=��'�9��j�M�n�`S/\������Y۴�3���aRX���7RѺ#���������)�sLH���n�3�Ȋum�V/�����v�́>m+��2���(��%�EG8G4K���xLB�&�y�� ��$�n?��*J�\YV�����]���W�N��$a�)��$S��Oc�e�&a���Z�ʖIEC��cE"囖���#��pK
��{O�Y��}Q�ss/ChF�E��1��:�с��Ji{w��o�x��gB3��(G=��g��2K�n�p�c��;`�UsqE�T>m�����o#S�rv1�t�)�i�K�E>���S�S	�����D_�IA�*8ԟ�P��Z?h ��	���3���[�
��F[�����(�K��ݭ��	�*����+^O	��/g#����P��2�A�h"7��F�?��wFu(�8�R�u�PU���9�]�����S��ͺ��1]#�=�Ύo��q6�v��}Y��يy���V�Ά3��}ǌ���
WFj����1O��W>n e,-����M�9��ܨg�&>�X����Х����^����_]��p�_lU�~�ɓ3���/�&a�*���lC�bԦ��`f/}"����z�~�M\?	��GT��	�%�R���?s�Β�Kz�1�}2���H!�3��5h��HV��D<����+���H�������{~Z�:�Fiu(��≿� �ӻ�4/?��2H�OW���Zu!��
��j4���ŲUz��s^���ъ6��� ʱ�+��U�<i�baR�ރXv0VPJx��AA��C����y0I�'x*�%�pw��i��)ME���B�W~��0-��3K��6�w�F�!8��EE��!�c'>�A��P9�ݠ[�H6.Nq��0�Y�v�Q��o-�GQ�0��&L0` �0O�4��JN%qR�O0�dVP��",�#�[i[%5Ͻ��/��?�� \�;�´+���3�'�T%%������Yď�C�G_<)
8�.S8#��'Qi��?G��zi��z��6.~
݁I?�V%�3�)1��ШU9��'���t�޼�a��Y���a����v�ԭ9g���Uwm��>%.����n]0���� #w����K�j���鹆ӹ���SmtrZ���}|6*.��y��_q�!���iD�w��r�Fp�� ^?n����b���5lVZ��@���$�I5Y��$.Ot�]��u�޶U��Y�$l(�^JpE�A�X��0TM�8þ�9�03����ջ�����Jd��y�J�L��$Bx�x2�Dv��[�����b�O>�p�B';�z�$׶�زe���ۻ,�x~0)�,l8���N�yeїq�W̓���f�W�"ErgQ��:�S��v�����M�~$��"��]�ݿ�	B5R1���x5�=Q�F[C������J��p�ӆs�NFQ�љI�_kt�S>鴨�-u�)�#j��E8�Y{a�?`��;=p���_��;�vD5 ���?9*�D6fe�ٙ�3���k���ͧ4�������F�K�'U)�˃!q�7CO��/.�6��7�Y�W2+�97=���7Hܰ,7,է�L&,�I믿%���g>Z�[�h�� j�C� �H���D>Ŵ�)d#�q�4X&�X�+2o�\^�Mb����w�9/����T��E� Ez��m��/��`�����^	�WX-� l�㲗����}�x��^�70���و��H9�WƢ��R��O-Q��|����Y-{�_��E���c1�_�	ݲ(ES�[������M���$jU�e(h�"
d~�E��ޱ�?�@�j�<��;�Z!���'x�߇���=2+T݂fФ.�?�W�ĕߏ�7�7$��1��h�}uH*��D˧V-[��@��v<�cG�;��JY��@��
�vF22�+a?U��Ĩ5�	%��'B,50\��Yٗ�������mcU����b�gA�}�eM�=�k��죭�w��c�$��m�a�
YH.�{�N��
K��9s��s1���Hq������R�oi�j�0zHE���O:�~v�x�%���CN�[{����ܩ�g����[�K%9,lX1XK�Sb#&
�d�k�����*��g%I�I�B��SZX���G'����F��uG��ѯ�N�X�o�=	@�Sњµ����S�X���g3�J��*	p��++�S�w����%O����骾?�a�!aE�l�q0 k��ך}*�� ����cꑯ�&��{�7k���}�+�ڍ�Z��G�F�X�3���-J�F�F����U���6W�>#_��a�C�=�0��#�×��>uU�����Q�o�5]��� N��˖'t�eo�rxC��t�D��?���ƹ�T��h�u�k��j�]���&W7���
���"��ddh���ϐ�-D���n�G��֚����]9��m?�iն�B��=X�PG$�LNг����O����P���ۆ��/B?3!q�,V�JǼ�ީ�2<�_^���!�n�6ݴ�}"�D,�Sr�蛮�]���{D��xa I<�(S�B$ջ��@?�q�ҁi����yA^�E�N�IR(c�4�Q�v�ǁyA|�E��T���}��U��'�b��J��'��5�\�S'�#�����A�~ g�+�c��k��I��IA_�c�6���G�!�K�o�w8��Y����]h��WB���&�O-�>�ϡ��"Û�^D7�(�+��c�"Q�B.�؂�����C{�!>���+�;DL��j�1���1�Y�
OsU1}ĳh@I�F/8����&�n[ǧ�t,���6��������;J�X�K$䰦�=������F���� ��&�XFբ�4uѭ� oq�'��l	�[��ʱ61�e�`�AϚ7cn��X��a��>��x�u\8���L��@
o�[5ѯij�N����Ϊ���z�W�1`�G M���)�'��t{�����;�R=Q<�2�W�!x�@\Q�rt���ٳ}���vMMuv`Z\�mˡ�
�t�䡮���<�&����Rl�����,׏M��D��L��I��I��ȍ/�G|�zNھ�@m�fh����c"%�T8Bv�4�a2�3�c�A1ay�����qnz�~*��UYQ�����yh��i#8$����;�_�����e�$�Tn�Z�Ax�d�wE�1Pc �����9�91e�O{�B&YHxQ���s
�F@�f�1�kk�,�b�k��i��[�J��x���g}�2��2=��/��,�2�@n�Q��l;;��sG����y��;��+ٟSo�1�
)��K}�5}���A�	��[�KFV_eiYA�A ���P�*�?������� �9�
X��Fv��Q�^�K�"��('��%̼��E+��	��@~��#�c����%����<r7�7g\f��!�(e�����u��7���i��� �k	�5��' #Kr_�igǘ�]���0��S��x���4�z�K�����vW� qn��L����� @x���RM~U-��^g?�׺����>�m�ûU���f]���p�xl�l�ۄ��'���xB�7�� Gb�X"��xR/�9+���əJ�\����"���D��%wBǝ ��?����}ٔ�L,'}����?��n�U5R�HQ��D�(̳FD6��x��-�ѫ���~�u:bip��{��7�����4��m����`��w�u&(e��j�JN���U�S�s9~��k\,Y ��S���i��a��>�3�V�i��/A<��]\'��AMyK%o��(� �:w��}Հ~�M@�L�\[Bi�~��-Et�K��ヲ��o�@�&�|��c�iA�`&9u�,[��@.��3���Ȧ��u	o�rQ��<䡌�`�CO.́���D%l	Ǫ�y�@�Vk����#�V�[`��%�����{L3;���'H%}�3������{������_�G�j)h7��t�8�,'��酪2���ᮟY��t�q.0ǧ�����1!�3�ĕ�oҨPk����������	��i�4QIޜ�H�U�O�Ϫ+gb�*T������'^	B��G]˵����Sw�F������d�Ӕ�+���m���\�|��뇷��T���1���9��70r&Q.��~�?����1���l�=m��_�t5���W�O��Ѣ����� T��C���i��E�"qX�}jT�P��yn��K�W�dl�������C�J���y�	�8�+�߫㱓��D�N�6PC��_�%h�k$�'�]�zB���d�eL.�rx�g��9�0$e�,�,��s��y�H�q4�p�|� f�<�"��(Q��-�t�1�.� &��@�YyV�S�
�]�]��d�d�wR�!>����=��[�Bt�=�6���Ыb�H�suo}Q�	�I��kO�>$����B�)��C�-�A��a�bS�Hp�.$_������5�i�;*�{�f�|Tk�3p��k	e�B����O�=DK�)�W!쾊C*H\ZV�ҹD���i��'0W�wo9R!�̀T�H��7g����q�r*X�M>u����Cw�k�CEQ���?�:�S��#�ԁOF�ӵBK������;�wCa!/W������A� ���C�m8o��ꯄ�Y����r�{�{��㍚'�EU}��w��B������U٣�����������C͂��l��A�O�*@��飄�|"{�4���U�E����^��_�W���^_�v^B�6s�(�c��U=��h�\�d����]ڱ ï��|��꿫�+��Z����'y��B�XY7TX���[�@���u��_P7�֊��kƃ��u�ړ�#����r-�~K@�f�<(^���+�eV4��|��忢v���2͘�a:�������l��,�ۨҴ5��W��Z�m^����
b��?��X/Mst�kv�w��֧�__}r �(�a��Yï,{�S<N�ٛ
�89n^���׏�N+�q�@�eA�-*eo�x���8hEꫩ���X:q{Hv�O%+�C)�T{��*� �b�����[bӋ9G�1ӭ�S�7&E���'��ï�Ѯg�[�I����w�X�SEGb�ԥDF�~h;��#"[�;N�Z��꾘�G:S���P��N~!�DkH3��:� 	�^+�������/����iQ�DS?zM!|pi��l0���(�r}��Z�T���L�&��ղDL�^+*�i�)�B�/��!�~6�H��
k�!x��(�֒`M��9M_�v���X��_��n"���xUNC�ͽ�o1��F��;%���;�q1@P��e
�x>yt*��?R���E�2Z3�CL����j��ə�q�7�N�Ń�=��d߸��������-�b��i�GX�t�H��x�[�Z	��D��}B�=�=�PB;L�В���љjm��bt�n���,C�B��3q�O���e�wh_�*#�<g�_�k�H��Jx�}!(��rR
9��wQ]:xe{+������(N?$0=���q,i�Q鋡0�^�M#(	IM5珊�16�����ِ�v�^����Uٸ&��wJd�<�
��5"�S���C���m b2����ke�I�ڐAډ�c�p16P�4�sb�!��o�v��w�>Yψ쎻wh�PfW}j��eL-�w���"~�S^_�g+���c7�A����}��U�)C�iA!YP�"�<;M�����,u��e�oO��1!0z�.=�@$4/sә�r�]i�U�CN���-6�6��	���;�y��Ux��X���RQ����qkwj���;��-�Ѩ�Ao\�'��	.ct�����/�q1Re+"�<ʝ�����x�!�c�	b���N5ۃu��È������ҋ��ʱ���Dj뼉,�Aʒz�5�,�.G[�hg��B Pt�%�qe��vp=�V����W������B�%���7�ݍ��8��M�W`�#\JĊ�\Vȩ��\�)�0��Ŗ��OR�E����b�+�J�޹_�-L>���$?���,m�h����c/H�X�56B� �m!)i���ÞoQ%1�8=��4�����\�Ty��.�z~�n�Ve*�PYLi��p>-�4f���u$����T����
���e�B��KKZwʉ�<�E9��c�'K����YN��"��n{�V&Y1�zQ�s�{F{��7L1��χ�E�&39i�C�����x�>�g�S�^>@=�c���H2��.nY|�;��s�o�Պ��̅t�b�S*�m1�)y��KX�I�ډ#�	������g_ ��A�xPԕ�4Pm��?�*��?2�����Z
V�F�;q���}92�K Ӿ���� �C�U�+���	���X�#�#�����Z�7z��l�7"`�#�ms(@���pu(L��*��2��l}P&NWͰ&�c=s#�C�`7�|i��,���Jy��F,ـ|��U�X���D��nչ�MhW���,��g�ĄM�- ���Ap�M$y�� �g��Q��`���W��C9Öl��Y�]M'xp�Rly��?� �Զ������&���bT�5����/3q��=�Bɴ�\5dH��L�ֲ%R����?)Y��8���g�[}(ǲ��W�ө�z5��IHLiXD�\�}ؑ��q��<�s}~�4�:��ik:r3�W���	74%\����ŉ��nu�y�x$j�����Up=�s�'�G�T��h ��Z�
���o�i��aH	���VƨV��"A7�d߸�~�y��yf!zW���]�w"���M;m��^�B$��~ɜv-�>/K_ ��g��W��;E���c�A�2�9��d[��{.���fm�#��0�o���Qˊ����`ֳGOi7#�,�%g/���G��V�)�c�#�qG[�p����п���\R;w ���l�s>3\���.�'$��汏�^�G�?=)8�^�$�8ٝ'�aׅEFM��h0��'��/'q.K0��wB�=�3Q8,�1�,�K���݉�Y�D�Eh�WA����"����Ǚg�l\^$��)�4J8�8�,94]f
E�ְ wkw���m�I��t'�o����m����O|�.(�B�9i���&���}���r�{ġ��8?$?��P}d�)�mlLA�����ךU5����8O*OƢ[=e���O�j�ڇF���QE+#X{��T���4m�f���u��m��(RJ�L�y��<��cϚ5����Dl3;�Ę�O����f�_'�F�z�-��.e�2ՃM7��z��z/0��,"Af�.ny��
q�,��Wn@f1B#"{��Q�#��	D����;�����4�Ç��&���]�������R�����=G�[�b��x�Dp�ˁ0I�7s0�Q�a�I���k*sW>_��c0n)�Eǈ��F�zaХN��h�p_��_9v�9�5H�ז��*Y�f�@*�\W3K��kVE��ݛ}�~ �wS�K:��)�s!g�)C����Tse����i�W���9m%��ۖH�~i7�Y~��9�z�t�uކ�7>��%�^�֍
C<���~��:NL��8�#LWYj��N���9��L�M��ɞKw�#I/���;�� �y8��m�I!��݄�\F������������h��*�\}'�n���"��%n�e�پ$��>��҉��� �N�1��IO5n�����
�|�k=������E,�m�Y/b_K�!���/�����8����C�U�R�hʶ�d4��Ӈ"����6\��Ŏ�fpRZW���	�p'����Tg�s��Tӷ�Zբ�{���d���O�7B���p�{ƞ��u>�K��HT��-�F�@�!f<�x!���5��sq�6=ڣ���v���2h�+a5A��z\���0�,+'F��/�).-���\mY�*An�bJ?�KM��kQԒ�#�'Rh�z{z������a�KY>Q�{�$!N�
��j9iE��)�׏	�q�	7�Q���o�oH�f�E�]�G�B:,�pv��z%��C>{1�8�P��]\m�8[{�9b�O1N0{S��Z&������X���g���I�����mXk�G��ݥ�e$y{�V��j<N����e׿�oDSG����I\�ğ�3_%��|�	fr�+�jO������B������?5�O!��ƴb7s0�F�c*�}`"N��L�mv_�M#&"��->���+e�����Š=U����h��c)ᅯ�KM�c�˒��=�4�_f>��d��s�F��"�I��0ӅU���͸�@o�����j�V����E�L[��ke��Hx91t�cK��ܜ��'¹�A�!��M$j4-����/75���Xu_dZ)#��w�yS-zEL�dNG��r���֓�����"�۸��=��sP=�L��T��B��z��I��g��Bu�^q�D!�2��E��<�⌸Fb ����}�G�f�rL�����]�{�Vj���9[(Ir�$��|����q"{>i9H�|�^����!�IHb?��V��썚�:�er�����-��ݳ@�U԰��wqJcu�%�5�7S���,��w=\ ]�����k P�I���AUR�c�H�6�h<���!�G����kw�}#Y7��	�}hd�.W�H�\A-�М�W��"9��^z��E+�"�cr���x/�x'V԰9C�x>!t6��^�;��=)���g���'dї���Ox��1<�ĩ1t@���/���ԋd�@��G��ZD�6��m�V���;�����������O׹���(�����mE_���PG�ȍ(ѣOo��'J@+	I��Q������Qe�2��7�\�7s҄>�<2����9۵~���u�=͈��I��4���k��q�D���d�| �z13��'��G��`�#C��]S�tȎ�L�^߱]!=��ֵ
�WD����	��cЕ��������s�M��q`��w\��g�HJ�����%���4�2M�R�ہ��"��'��z�&L�+��������P���$/� 5��=��mm����*A��ܠ%�#688��4\������w��y�G�U[�n��*�pYG�o�����ё��{$yjƠ�܊��|�� ��e〗
IZ2s�����E��ic�Z&�G,���'|+��{C��YL~�Q|�os�|�F�b���1�� ��ɇ��&i��~�@/x}�	g�'��i�=��x	�2|A�n� � �;��s�}�%��������9S�?1)Y�)��`K3����z�$%�	��5��y_��A�(��PH
?�2�ڞ�Ө���<
�@�F�}���;�g�K;���^�+��w��`+�PG	�t)W#���Y�K����2�(�A7�`�>(���8�(yRG��u����֋��n�	�'	AQ��+�<�>sV#�4_��x��w����g�Aa��4���-��0��7ȝ�N�M��D�WW���O�z����� �o��|wM�����g�ʫ��2��ݦ7�c��q���Nk�]耂pۦ�lf����Z��e"��}�ӻ�R�;�b��ᑢ�/��i��3���^�\�A~�ؚ=Ǻ��%����J?����T�΂X}��?��������59g�HGW�DMcM���ޑ�8C�#��N`�~sU:���if�>����¡$m�4�{�Ñ՟ �l��ސu�|Bjeg�/8?U�Fs�����'��ð �>�<9]��i�i�E�a�]����V�I+nA2��ﵗ4+�y�=���i���wN��ն�]M6RP�D�B��1~�e-;)�K:�m�(�g��-��6�W�2�McX��A�$�9kI[���.�����W�;�b
9o^��Q�g��m`�C�O����º%buM�`�ua�V���.�#��^[֗n�[>�к��1��;2<n��37y������፟���G��)S����T8�.�'y��y$����)��x4.f��������x^3��g�̌ߨF/��8;c���/�.��8@����嵚��i���gI��ő�*D�����Eg�g5]_�Ѹ�w�~:�|`_3�B�Zz�J�CJ|�mE�&����|Ga�����T�������(�?r\�2���p?�����D��l�dy�� ���C&5*jx�	�O��:��j���� $���-�� E�C�Xv�2T^��������Z���gV؎F,�J5شy��4�[�U���u\D�7���W��K^n[�Åa�x'LPz�b����eB��(v��ݔO��0o�,}u͛�-ay��q*�]�2X�flgp"xtQ����d����i�VJ�����a���v�R�]������Rb�!��|N=�[���P?����w��� s�Q�٣IrYk^>�'��=>)�������a�R�>/hp::e_O����5�v���*I f�� Jn�3&�nk����x��yw��҉�K�̴)8�!�WC��9�O���&��j��Wcq9�I��v��Hm�7��ו�Zu���j���%>��������;Cw��m�5��	�1#�T��}��u�Ր����蛊��!�w��/�-�	��2 ��psJkmnD^��+a��S ڏ���h��q���C �eb�}�Z^�����H^�� 0^��߭ѹ4��w��Sv��c���O��F?][�ٰ@|��+�ꗝ��5E�s�T�_�Td�Y���`9�J��$�Z�Us�Yh�0nd�l+�B~�6�ȩ�[ˠ}[��:�Z򱞉�Y'/�"߸ĵ���TN��5ou��^(᝕�_�7���+¯ƹ*�u��i���$�X��-,.}@���<޲�l����v������v�{I2pa0�X��x��:�(�K@�,�R����>�d$���\+mTH���sb�Ȟ�^�MiA,k,>�^�;�,u��5����a��Y��{��NU�M
@�9dL�ׄ�ߏ�n
q��^��A�o�u��E�/���:��|v�%!;�C�J{l ;ݵ��X���G�[�Be9}I�1�ҺS�׎&��>�<����;�gV��Iݷm�m��XFm(G��z�t�W��(��G�Ne�������S����@*�DZG���)3�G���	��\+�]u�(��e���۶��?���!�&,���0��=���}��Y�\ȗȉM����&=gDըW��\�
+�]��_���8r��i�{dr��~j�� ��?�֞C����4�/6�_����������U�}$@/�kM�U��ͳ�>o璒¼���q3�x���'��ƣie@�x4��t�"�㵇��*<�(�����ޅj��8��g67���;�g�sb�dչ����A�-Hߥ_�G�К�f�֮a�P�v��U���n�=)�@P8'5L_1ѻfܙ���X���$x����yB]�q��g�|���L�`_e<]T�!��p���}o�=��rȭ���]0�"{բ�)W�9(D�K$���q��q=��i�@�W��^0�iY;�IC���ECg����UfD�9����d���N�U����s��J�e҆@D5��S�#ȋg��-_ X��tLk�ݱI�DwA�:�c�@[6�[����!��޿,WGwi�lYRy�ph?vgW�F;���--�I"ϲ'�"�&_^�(;D�+�p�c����`U�sk����CM��!�<^(`;���d���*]�"s��_O3@�1W�K�$F�@�-/��I���_����`���6��{�����!�;��Y�	��E��!Ǚ)�C~��g�� Y~�	��cj�ў��o_:'��	d�M�̜�}Y���eaz��2 �H�U�?$�Wπ���ې�Q�uu-���a�Q���HM�� ��ɿ;�r_���Vaz�P��"s�G����>5�x�Vt|��'����f="Hȵ�W���q����:�x���[~MF}�`�.\ 1��Y���?%���́s�mĸR=uȁ�%������U���L4�Y��l��� �۫��a/����e�8>�m��|z�j%gX83nK4�W��dW����4y�;�0X.n+g�*�o�YBo��&����ב��I$�S����� ���me��aefZ�;ٖ���E/|�c��q�������wT�v-{�ݲYgI�Q���s�z�F�֓7�1���=�쇜иi�L����xXpg.��Ŕ�J=����ӧ�27�Wn:5DO�;�:6s��7��X���yo�<�US���1D�/)o�fK����BڿF�	�']�\Ë_��>AG�ԋ3�P#�d?T��u+����J?
�K�F����v��^Kv�p�����vg�\M+J��	)[$��#����}\�PS��-�2�77���Y`@�ct!(�#G��u^ǯ����R���]\tͦ_���#�E=�:�_�r�*��2~��)�C��v������r䪊����[�W���S��s��C� ��﷞MO!�ݤwgP��Dx������U�L������]��p�Syl��۵2޹
5.�0/Ӗ܎�Xx?b��%����/�?9糖����\+?`سG_��F-%H�_��S�?�}���B}Ν�}8����I�2�5�!aHBeZD�0��wNI�����CЫ)cR~F�s:3�ia�m(�����?�4���?��;<��Ho(u�pv� j ��J�Ufpls�(����C-�0 ����ʋA� i��a>�'��śV<���A-�(�nh͗�ϴy�y������:w�s�Q�_M1W���B��~���-�3[KVK�cr��jx�1�Z􍎪ci�A7�9�s�[g��.:2�ꜜ�9���1o��Qe���`��O�mb�b�9%]ۮǻ�SWV��89#h�[N����еC�̌�;�.A����3b@j��]�k�܉ˏq�GK��)nB&���8��-'=�΅{�3����jT\��.�b0�m�!����3��w�gK�A���ϧ��JM]�MPA���M�Z�&Ԫ��a�gsE��M��*�������I]�����w!���7sNN��կx�%V�t]mఅ���|��"�0^�o��������c��r�0y��X�?���Ʈ��_3FlB�����R�5�?��CO�/�ф��"B|�E�髐#��J�Ea�{Xq�T�j�ê�-���p�՘ĻB_ю�P�JЃy�iI������vDb\�����������\��'�yzs�۶��Ie��g����$�]80$,��4���y�m�q����b�f���"�d�Q���":�bԸ�qM��Ø�7/�>��.��]�I��u+�R�y��)�==o/[~�����z�p��`�his��{QrwI}�k�h>Ս]��k)���>�_�Ȋa�]���p�]_�� �o�5�'�L-�*�ߋf���ş�3D�k�$��!�t�&�-��K��\)Sp�!]�LC�a�WҊ0@�J+��KW"9�����J�HH�f7^%���Zp��+@�>���T��1}C��]�����0�C�dǶ#¼t� ��Dn����H?骃Kٿ��wTY/�l�H���1� �d����m	_s�ۙ����J�k�X���y��ca� �}]�E���֌����ۓ(�����4s���Ǝ?���T���RO�T:�K���v"|y^F��P	�KrEbg��O��_g�l�����S���p<��U�h��Gd�E8��&�Q7q�,{��{����$�Z����]�'��4�sT����T�l��)X��SB�}�ˏ 7�4�����Ԝ�u4@3�\�$˓��-�5*@��E<9��'�b��D�, �v�}v2�2���a+��0�����f��,!��c�뗟:A�+:�mO�s��hb��S�鑽M��Tk�y�������p����Y?a#�-Y4�"{y&�N��4
���9_s/�ߊ��@�q+����)���QoU�v͜4�E�!���:�1mv�
%��@C���{�B1�PC��S���[�*�9�(g1D��S���&�"�פ��H���mgTHI������1X!*bGw���o�����E
N+J�[hruIS�g��!�?x��U�*3�d�p	\��+�p�c�N� <����U�?���!ͱ��X��0��:��s}�C}�
`�#���}j(&X�,�#���7a�+��O���Š3�S��:������{���S����2�1Q��*��_1�M����#��Сv��A���fU��ͮ�oBGO�w8��j������@I|e�x/�6t;�pR��&L^��*b��*!�W�jj|��~�7����$�юodPj��y�&�|��-�jJ�Z�Gi��yGF��Y�˛�����.5�=ĆP3h�L��0���'�������\���s��V�B�U�q�l�:xǨ칩{-q<��k���ߧZL�I��}F;��r�/��C�]��s{�s�d>��p(?�\$A��,��qX��ihJ�2^k��tI>�O�b�}�p��h�ސ�\�@����iU� �����J��S�[��5��S��������< S�6��h	k��I��AKC&cmXh6oH�DrM!��࿇�w$�Ym_���UNh9W.e����-�����"��^�c����+~�vc��Ů���n�r�f��C�$!�bM�4;��/��ʝ�W��9�v��O�$1r!ğz@���/$1`�C�Z�*�T�����\6���z5q��;6�읷���
������}�^e���j��rf�D�	��f<љO�om�'�z	y6�G��X("�e���-{��x��)_r�;�z#��k>`�e�u��h��$V�����2�J�:�[�MzR���vzg�G�dGl�t��ZA�Y�t����WP�'@@=��ѵ	bJW�N�,7���?͕�DZ�n�,����M�M`��\[�bˍ����u��eè����[�R����w�sj�{�繰;QL��Mȵ3��5�g�����/Yy�f���S}�m�0��y���O|%�x8.Vc4?ţ*R��!y�~�u�nfQ*Q/lY="���E�e"�շ�$o���pL�K�H�V��e�\���Z�$����E�3c� -����*��r���n�{�Q?Y�4�QrTsv�QF,�Y�؆1��FϘ"��W��ifB�6/dx39�gih��/!$=͠��.f�2�4�nU���ɳ;���s3���[/�#w䗾RS[��1_�)��K�u����Z��	}� ��ם_Q(�A7�q���P���?�ڦ���3���Xa
DvaF�a���X�0�K����Ņ���f�z+��	D�Uj*I#d#��Ϙ������(�K��H7St�����Z(����u��r�̭�$�❀*w�q�!����>�#7w���	�mM�=���w�0q����'�溟έ l��Y�ܒ�W�3]5�񸌁��,� �����M�Om�ئQg�- ������/�Yz�'q_���]��p� �l^��p*ӹ%$±�A�q�ڦ��b%���/D�(�n~��\�\�؎��0��%�@X�춚?:@k�iP�θ��}����b_�Z��5o��H=��DO�2��"y������ ~�O:�b�i\Ř�;��١Z�s4����yϟvŕ���uv��^j�E�e$U��s�����/I��� �<��������i'�a�f����>Vw&�A(1���ŗ���y����[�lj�w��W���M,|D�o�MBUd�~�-1^CK��8��'��(ǫ�,����}'c�C�A4i9a�[B�L.u��7d�����io�[�Q�,�Α`g��O9 ���%Xa��8��CV����%o#C��[L$Ƚ�YFа����M�;��I4�3�{K������ץ�oG�)� Ƽ�:_8j�='x�؅A{�����O�`|.�+��觘��P73�[�*M�<sǤ�����1�e��ȇ��,�ވ���dɻ��g�a�@�x�H��qu���� s]7�\��(0w|���ai���P}#� ����m{М���|�%��s�iɊh1��Ә�Z�,���r�����6t?5�����U�z��l�6臦��K��5`5B�;�O;H���X�=�D��=��k���({E��YXl�kT^��e)E��t�P�.��z����JkO�y�E�����˒:���Dݠ����y��ܚ� ��W��'�	z.,���e8�S��SM�S)2���0��,3>��_	y�d�q \{��`f�G"Lq Q�����_����ɜ��-�?����!�]��Q���Rظ����=��'[Y���)'������Z^sa2CQ)*3I���k���>-�4��)��Ǚ�iw��a!/q�4lp���_Ō��
ѿ5L�קx�*���f�%@�3���k�vͮ���o��܈V�Kk0�)n�x!�p�C�7XF34�%����Ο �-W��%9��\�l2�H#��7Sg�S��k�e���D]>�(���M�g��C�yߥOcH�+�)���[#}���:V���Wy����>ٺ��w�*A/Cڠc�5���� ^<P��<m��`��'��m����[�h��g�����T��+}��%��M���.��w���ѯє�c����(��e��OF���Z��],|����)%�f�E��%�J�_\�)��9���P�HR���$����U��3h��}dE?%Ӹ0��l󁩧���V�˞/Z(5���'��F�._��5�TD����K�,i�^:'���H7S�ފ����.�u���7wU�η>-b]�@�P<��I��_�ъف�>E�Q�fvm�29#�a&�����f��nu���,�	�>`��p���7�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�+ڜ4X{^�wLРr�A�}���Jdq��B�Ϥ!>m�gخ���T����r�2����,����.��km�EZ2�X�?C��>T�Gt�U�����Z_4�ӫ;�T���u!U�Gip�L��C��S��S��!
,/�0
Tf���3�^C�Q�$�Ť�^��!9]�f`ay�ȳkrMX�6Q.��� �1�F�j���xߖ��0�Q�:��澀��MN2�x�^/hĔZԙ^�F���[�J`�&�/�]F��M8^q�-�Q�H����2��:Y}�Ц�����л��8"�b��G��Z�*y�p�]����*b2yso�Ũn�U7w�-��h=*�a����<Wr�ۤ�f�{�����w�i�|N� �y��ZQu����]o)GK�Oz�::��S?SۻQԼb�a��#�fϢZ2+�jK,%��p>Ïi1���$��28Rc�"�	�+�*�ӻI��VQ�X_��G���F[�Ow�Z>$+�����@l�W1���d_Dh&d��뱛�+�wV9�K����l3mY�p���3�'��^�'�>9x�F~�
.�B�U{B�g��b�᫾���f�P� ����q�C'N��le(?$j�����.
ͺ i�?E��4�����/zN_[ �5�$����ɿ��˾5m��(:AH$�pz�׷ߘ-���+��-�Ȕ��Ŋ6ǝZ3�Y��>X8��~`b5	l���yX�%f�t�E��,.�:���ꎡ-����\�s�9����{k|���.�M]O[�@��_�1D�B��)vP�{T�/ ��"�"�H����Uo<�<'���L������OyX��A�_�`XU�I���'?�&�W�/
o��2����G�{*�e@����<��]�/gnY4P����8�h��	�F��{%<2V �|y�t�8�t�ȖE���L�	S_ON��3���nZ������;z�#�{O㉨�s��U���IL~�j2P����h�.�5�'����d���X����ê�We���kJ���+1��o�(�j;��d�N%l�[�����J�*����\+�Y��x�׾�Ů�l��C7������(	�pqijc2z٤�'I�6�[#â�`!o_c�[q�m�����C����z3EK��L�G����ֆ�'/�L�X�x�η�K�(�г� ����\#��%�+f��X7��}%�~�0�$I� +�x]e�qi%�r�dC��]����v��m��m&����
�`�2c߉�� -��&�Iz+� �Q�X��>�ن'|�Du	�c��Ξ'�f}���f�( �[����������0*gB³���`��f��#K�Րx�q����N�a��6�(28B�k�ܯ��M!��1!�s�O��s����Rz�?�*���WZ�!���z��R��[_��^'�(gNv����ԳRZ��,��1�2t��Z�W0�gc�Tl�[㹜���d*AM=�txdL�P�)���ah��J/�תAcG1�ΐR��j���:q�iwN��s����b��$�( ����,�@͠@�mm���,$�����6f:�(F�6M$�3̹'i�o/dcBz���9m����<gl�;#o��)P�+h�o��b��3�1ܵ���S���싑ԉf�! ^�`��/��j)��o)8�n�5n�h�MNPu6S����筩HR��`�X{�*>��Zy���z����6���u�H0R�g�lk��&�1�\��;gS�����G����]�y̞�	d�����U "]1�g1�ꒄ	��sB]Ee�"�jA/��4.��H7�6�
��zrO�@�� 
�&	�D5Te�7�7榀<�����꓉7��C��D׃=��[��{�w�\�.g��rQ�F�Vcw�)�aḅ�C���d�����VG�mY�ω[y���z������Cp�Y�=��P���ſ�I�Б�[��ۊ���-kR&��3�8��R�ꊮq<��͐��] ��: ��QR�U���q�d��qɷ!�$�.͜�O���Fj��v� 0�ܑy\��:�B��3Q��>���k�z�g��ycľ�խ�K�K�x@3S�uqTZ������ÏZN7�q�`��SU��S���f4��h�dmS�-U�
n�.p`����3�����Qdt��)'�Ci.-�'�� �R���� t�
��Tl��f"�g���!k������5�#)!�M��YJ3��pc᩶�����x��������;���'n5���{$�k�&�;ų�22���v	T�0��na��S�[*�8�;��O0ȽkiY@&���@�sJ>_�e���Z�]֏�!ȣͅ��7Zy���
�"�� $�?���_Zs5Pg:
f�%4o�	��e�x"=E���I�4Ѭ��]4|S�����Kor��t�+����) ���Ig,�
3{|�S	!`&,�w�'��`Ц7^9�I>�ێ
�O��!�D#���$w���t�ڻ�1���/锞0EXG�ͽ:#��tu9?�4�����zQ>�1�0��U|/�b�!!uq��?vkt�F��C�}2�ϑ�:�1�צ��XdmI�����U;Pn�@ү��+!�ܩ��)A?/h������rk^��CW�t8va�U���>��5�f���S�B��ݑ�ǽ�K��Հ�-գ>��I#��P�tXo��ܘ<:O9��>�,Fgݤ�K��G5e�b��DI��U��Hqz*���������gH�4�]e�A*�]7Y�6�{�?����Xq�C��Wŏ�̮5��\aLBcmn��?U��D ���d1��\2�2���W��Ll�o��se�rڽ4�����Fnٙb^�1��F�:j�u�MH�SLZ��Mϋch��0��׭խ ��>�C���xu�E��m���
4G� B�q%�w������3�Z�͝;e�_�%���_���
�L��3�(�CZ��ο�k�l�����aך�z ��������@�8]4ہ?�B�s��Y��F��%�F�IRo�֣��&Jơ]�S689�f�[|�n\��KO���3� ��?8�h{^�	ˊ�[E[��� a��eKl��-5Ў�v��h���1�����Y�1��=���5���<x8A�_��y�����
E'fC�Ԇ֍s�{��d=�������a���͡j���<�=���Qώ���.���vn�l�B�3��.� ���=�:����U���kv"��[t��[�!�24�����q�U���iH⊓���ϒ���ޛ�5�0[�Mbh)�گ�*nѬ\O��Ufbq)oO�n��JwL�s���*��܏^�e<����y�����5��^�wq��|�]��n8��#Q��\�����Z)&�G}h������r�?�(�Q	�j�6��#eHآo)W+�},g�j�e���$|��'���j8z؜٣D@+8Pt�@��}�b�<h�u�`�F�ұ8Ч]��ʁ k)!�@���3s���~�A3����B���M`��,��U���d�$&C�x`�_�E@[�Z:���1R`=p�>_�Ez�B��)j8�~lj]��-F�[�� +P�N��(-�����
��ړX;�M�F�+EĝXFsww� ���A�����D=��M�p��m�记l��y���2�\���d�K�ۆ�m{�V2�� ?��>��TG���Ȋ����Q _����&�.�yT?F�uk�G�C�L@V��%�ؾ�9!լE�[�T����YL����Ү�Q����!yf��@�S�%r8�Y��Za����<sa��7���XU��Iv9��<���
`�M�YMY�X���E���=_q�-C���i���]�b�CaC�����n,�5U��P� �� �0�qb�s����t<�s1S\��߼�H.a�}n��6��i(�@�	��nJF���(�aC�N��-�S/|��w���)��]�Q[s�N�D̝c{-dj;�����v�(�w	G|J�p@�M1%clB���쾵Բbt��.=;B�~��pN.z�U�n�a��"�[:U���=ư��&[�տ򝐘���#So/�R��Z{��*$NQE�D}�ZQ�ui�ݨ����(H���U$��4��?ƶ,aT�)[V~����i��Z�6�/�*�B�>2�$=P̠>`~Ӊ�cF!��npg��R�ط�y���]�uPT����)�E�����tحP �k�"jGWAɚ�2/����\��&j���wT��vI]��,^  ,2ߗۗ��FD70��ǌ}�~�O[`���s��?f���Y�|�ku����1�3���i��a�"�<Gb��Y�	R��+�5���a3�@h4G�x�FQ��&���[�]A�@�pf�i�<3�������D�_v�+N>�@}x�e(��Ґ��1���r�X{��tѶ=������P�����L�hdF�
�^�`((��Z�K؊��<����y���C�9S�x �&�j
ق���n���P+����eN1��ʱS�9b�u��q��
>6��%Ԝ]3aN*�3w8`�m�K�~��H4I��ś�ѩ �`���.�*�wu��K�-˨�E\�TZ�:J�N���&N5��o�u�� :�<G3��FxXO��=�2����^gi[0������\,�?}��GO�jTpE�����)�)hq��O�9\fܤ5�8�0�ʹ탶����x�)4n��P�z�
{ዲ�d�}xě7�KȆ���������b+��$�F�U"/-��H�p<os�lX�5��sG�N
@jIzKY ݛ��S�����J����8qQ-j����)Z|w�e��ī�b+��ü��	ʯ�Hq}���QmRj��͍Hi��RV\m5ò�e1;뺩�t��	ۖc�b8���k��l��,A�h}�0�PfO�=�x�D���k������%��o�|�=ME�!ˆA�7x�PY���{
Źi;h���E�Y�E��
�б��{ jV��v�,�17�3`�l�,�o=,��M�y{f-$-7�q-C!�A}���K���7,�tF�Mf�cV��A� ������9��>|�z�_��J�^?��\�@V5�t�k�v�q��
ˣ��R�fӤ�QXB�%��	�s���+�����@z�Rr�v�J;�:���ʃ��&t�r�UkI<�~ߙ��
��>�
:���"�L�c&끲h��(U�/��?�3g�� t��Ja �y"�;�059���&%B0[m�k��O�1�aoⅦ^�:3�_R��%;�o<VX�����X �=�VH�@�EE�A���m��a���*~������6�i:�˟6L�9��yG���\:�'X��7Ԅ�+�����z7�a�L�"�H6���*9z�~&�($��c�IO��ag�:�V�3��P����;�	�<�O��m�O$ �Wt�uH������;.)X���U�lQ�LdSq)�qV.�H��m^�,ڇ6�9��_�K1���i��ڑo��(���a_�c�!p��a�k��@����oS�����qe��Z����A<"�*>�ɵ)k�Q��������NXm��V�.ʷ\]��O��7�&��`󪣞�ߤU��V#�;�9�h����_�3�*Q�S��/<�('��g*q��K}��k�P�񰁽Tպ��BqHD��*C
/�~��3]}i)/B��O�MiN��W56���Y(
7	_o�8�V���d,��	�W:��\�Fϩ�=~�Jл1���+Y�d��J	3���TjR�*�ue�91"��vkB�6���\Q(�de��}Y������y�<$+���p{��`$��Ѩ]�0��%�:�&��a[�=�${��ۥ	�)�r���S����6t���G豶��d�v��@1Prr	}�Ô��S�#Q�̰+����cK��TלPۍ���o5Zv���Zq�j_^�=���&6us��xꙧeޝ��k����Ȃ-s!�t2�<&������83�W�w����
!��es�6N��cŮ���n�M�r���*��A��1z���q|w��E�s���Mtf��0��ܝ'(�/�~+���?�����#&�4�OU��9'���,�My�������V�0�!4b�}٫�2Ƃ�R�A������ŏ����F@PӤ~KR�'1ۊB,������s��N�\���V��ik���5��]c`Ru�-�E|��z��4��W%;�oG�p�,z���ⴛByw�#����!�#z[l��&��]���I�K^O�B9���dV�TUI��eH��_{��5D��B���l�� L%i��*[Y8���nA�F.t|�`�L���W��i=��R:�;������Cd�D��t��>��U��:'Qd�P���6C�v"�@�i���dT��l��^:wOP��iu���v��A��q��w��|?�+�%��=���a����&x �Ě7]P#�Z�S[�9_D%"���ϳ��&Iӯ�, ����������x����� u��^����d��c.�;��� "�K����ѬE:^�)C��apg�Z��U/�h3�Yb���� 
0��F���߼f�G�y�ƌ�и>I�ΕJ����}B0dh�G}�̠QJ`~W�)V�6b_�7�J�n�lwŅ�$�d}�:ӟl�`p�~ׄ_i>Kd�h�� ���|�(9V�����l�q)K���������ã�'y9~��3�x��
g�|,v�ǲ��hؔ����n� �g!�v�Vh�X�m�pe|�S$o�D��.O�! NB�E顲2��I�z���[���ɑĲ
(O��O�����M��H�?Sz+��ߝ�����.+�{vԭ�J���.��d�T�X=�Y�#{ebz<��B�y���f��E[/ .�@��ǽ����O�)Fs����v��{��J|�A�.��xTc�@2� _�N��'Q5)���{y� �5�͇��`U9���d��`'����Ly܄`�FG�ex8U7�r%��'$�&D//�b�����%G�"��
����; <���]���/�@$4���� �m��	a��dl�<pK�бΙ���9�f�����]*	���N�����Z��)�Z�H<��~<�{T)ɨ?z�ǚ���.�������hZ$�5ւ��jS�	��#�|�D=^9ނ|�k�r�RJ
�+6������s������O뗀p+vݡJR	���!\�D!�A����A��3����{�=�J?�(�^q�2�õ����I�g�6����l���#�_h�1q����>�(CqZ��|K3C�L���M���Z��ٻ/��X���S� K��b�xR�����\(��%o�f6X��}����U�IyɊ����vW%b���ƌ�B������A��dq���-t��c$�7���-P���nHlR��Q�Cj��(�+����I֪���bߞLܑ}F:CfQ���`0�ْ���~�p*��+��-{�%@�f��<K���x��%�_�Q���ca(�ݳM��8`�J�&��Dm�D	�θ�u���R�fצR��G���!���&�n�TuR5_���^���gs�"����9��_�<,����vH*t�}I�܋�g�~�l����fB���A�tz�h�t]�)aaN�S�t�>�L��/ɢ)As��1��y|�H�����<����'�������i+(�d�l������m��,)�����6���(+�M�Sr�X��KV����cG��L�c�����!O���8�&P�E���n��g�����Q39��ܚ�%��c��V�Nu!�EP`��Ω�B~jn�N�T;Y��yn��_MT�6��f���N��{X�V`{�Q1�^у�FӄD6,1 ���H�P�g�?{��b�1!�`0�t�Z�P�s�ьg]?M/�R!��
w�/�P"�O/�,����G��H]�w"9(Q/�U<.E�<7&0��ϑ���B{O����E�!�k;�D�eE+7o�<u���x�Z�� $�҈+�D�V�G�֠��!�잓
_��HCn�V����/�bQ�븵8��W��w|����VD���D�㬸�E�����pR�=�����i��d������)/<���k��XR��/3�.��p���×���9�s���� ~}�R[��Ȍgd;L�~�	�)�!.l�ti����ۼ�0�,Uy��:����!�Q��>����߅�g��y�p���Kα���IS��WT]#�(�}4�T�7)�J`�y���S3�-ؠ�ߥ�drB-���n"�`��^���0�$�Q)�c��^��H�H-u����3�7q��>�8ň��t�F35!��̠Ck ��i65n`nN�e�Y��>� ���N=���ӹ@�+���q��!n���>d�=�&����y2�ǻ�w���ǆn�=�S�S�����\Ȣ!�i޲��ą�@_���-��j�]������FHȈ�|�Z�Ϲ�	%"j�)2�bc�Z�,cg�fr�o�v��*�"��1���[4v$�Ӣ��|8���*F�o��pt�2y��e ���Iy~
x�U|�]@!�lD�/��� ��Dj7c:�I��M�O�'�����#�
�$<�������B�j�g.`�0*�W�RnQ#Ư����u���4�eQ�tFT>�q�0�'�U��*�!�OΊ�rn8�-��1��I�g��#c{�s=$,�E�����ݞiz�@�-���d����$����um"��B6�Ght~u�������Z6�{����B_*9˂�4̾��~�8c䫬��N����ؕ�]y3�˻h�P8�?����Ҭ��Q���؋<��	+j��ɸ�2y��Y�qa�j��Hw2�,v�7� $%�2�@חf��D��t�o{�[����2���
��Tc��>��Y;S��%���1z�[����� jzG �Y"^��p�+��V�K�3��Q4ep��$�E�������]_ �@}R���63WB�Ɨ�����D�jK��N8�s@[Xe��U����1/�ɚP>�{Fe*/�������"ދ���B�h��Ě�&���`��:��K�bb���<D*��B����^91|x��	������}�L�b��@���<e4�BN��x�hf�����Z`�O�1���l��{fPN��3��`42i����ILVb��� �����0$�� u���*�A�����H:�$���h�f^�u\�d:�J�G��F��pO�_W�P�K�Z�g�P/����T\
��}8��Oa'gT�pD����ஓ#)�/l�m��\D�v�OD�p���V��gWyA��)}@ln%���.xHztR�?�M�[��˔��l�������ɱ 1
0�{�3+�U �Xq����@m��J  5�����~Sl-9j'5K�����X��8�ܯ��=�$�g��v78��.j�{0�J8|���uĉ�夡D�ZM��U�	�2H\s�3�R��]īOFi'�Vp�5ᏺC���WA�ҿ��'�c~"Q�F�kC*l� {���0"��Oη�x�ו%/Ykኪ�D����B|�VE�M��_i�xi���;
k��i2�Һ>���r5EI
������?w���=K �
*57h������I�,y�fM�-C�T�$KJWq����S���*,�*���ץ���&�_H|��z��A)S����>�8U�=r�J]���A�.�^��Rk�o�ϊ��(���z���9��X`�%�nI���fG��}i��rt��hFa:�9`h�o���r�/'��~}!�h�\#:����!�L0�F�Z������̰�����Q���ޭ ��a^��""����29 ��&��N p�IPJOj��a��^�|�63mӲyɩ;��<5Y�����Ӷ23 �_��H���W;�De�4�RޒL
}d�D�VT3H��mH��W9*��1���H5'rU9ڷ`\����Q4�����p��y�Q������S"����N���G���0A"A��9����w:��� =��mՎ�LIm���Vu�շ���r���!ϛ�y����{�V	T;7��hz+�-��/Q2>��{�(MKv�M��r7}n�v��gq�`�iB׍o�%�
��G�}ϱ�B�H�Of��N�HoW��.��
�o��K�(�c�d�������W��g\��^�Հ���o#1I�g�Qzbd�;�	�}�U���z�������1�[�v�)��l��r� �2o$���ݣ'���wFM���kK��
����롮]�IK�����&	[�G3c=-���0E�	��%rh۳SY�7��W�<I�-F2�J����@WhMrX�%�i�ۄ #w�
̖4�R_������7f�=�P��Й�'�Z����@,�q](^gc�=��r&b���R�ʽ��hok��"�no�s��qtXQ�&����8���W��ɀx�!ks轑����Ŕ����M?=�Bo�����i����q��/�+����M�6o'oNez�o��'�/q�5~����?��
�%�#�I�4��U_��'c�O,��9y�;�����i�V�4Hr��QA��H*�g:鎗���k���Ff|ӊ��RK��������B͎��sXq�����|��OS�/��9	i`x��-�b��K�\�#��}�q�Ug���z3����gB_0#*�;����z��ˇ��~�����B�9�
�mT�C��E�E�ͽ�슏l��J�Ᏸ� ��iq��*�f����dA���.�?����&gW�STihC
�xK;��r��EC�ͽD����٧ۘm�G�'w�-P����c�FC�EB�fb���յTt]�:2�^`֖P��u2�8�ܳA� ��֋:ó��W�K3D�#Ð���@��xBhq����:�����[>��E[^%� 2�尡��*�I����:��^�#����~?���'�;��u��^�l���e;�=����=��8�"T$w��1�k�t^��:CIU�p�$��y�N�Yͫ,�0�����������
�ƲÀ�$��ݾ2SJ���%��O6��2�EJ���W��V|��_B7g�p|V��Qwkz$6���`bMl��ύ$��_�CWd�8���"��9����%�l��aρ�����2Ʃ h'Œt9�b2~�w�3���{͝�R�ƭ� �i�/������OD vm��y:�����Oebc$����L�.uH� 4�E��زO���z��U[���/�ز0�￢a��`j*ǳ�MH�zIw�C�X��7+�ԓ����7�(XS�D��:)TX�$O���	b�5O��`ay�օfN�E�KV.����m{��8`5�O��s�t���\{���|�#�.���f�@�l�_��{)�99{�� �� �m�⌍`�Uz����ڭ'�y/ky�F�y��sU���K��'
A�&�6�/�3ǰ���ݡG����p0[��7<��]-��/�t4;��������N	�3�ʊ	I<����ND��I��_^���P�����	^'�N"p�ǚ�Z)����t�n��d��{�Ш������!��/���3�`'�h�p�5��uX��o���I�v�u�������[J�:�+��}�z(h�Քe��Uގy�������J8���DD�\6�:�g.��!��ٲ7�+�Y�����0��(��Cqty�2�ɤ�I<��6!�������m_�q�W"�d�eCWF�¥�K���L�0�g���j�u#��/�yX�6���dUKR{-ОB՝ԼC\�+1%��,f\��X��}P���3RI��Ù��/P%ȉ�����(@������u,���ò��_mKV�k��cJ����-�g(���`�>��9�o���\�zUy�@oϑa��~�f2]E�F,hn���C�����_��x*
�d�/�� �F���+��X�h|w�P���?A��9���� /��_٤�0{mt���S���G��ͣ%2�C������L���<�m�S6*��깴M��;�"���Ι�/��t�6����	(&c��$N�5>��F�m�Al,
Qj����6��(lW�M�����w�����c({1�MW����b���!'pϕ1KP2����^�H����}�3Z
_��{�9T�ϒR���g!Ff`p0���j���ܕ�J�Tĝn@uM�� 6yN��zǩ�A����"{ �D�u�M�p%�c0/6�@��OHևgWn��]1�x����YV��甲�Q]@�^�.�E��0���?"���긤�˸��]�&K"Za�/��z.��F7����ps>�X8O��;�F({��VD[��e��7��<��9�-���\%��ҩ�DD�� 騏�!�K���6�T����)"DڒV���O�|b�]��9:(�Y�7�� _�Ǔ;�3t��ip�$�S�����[�p�*�=�����{�e@�K�:����k����B�RL��3��e��/A��_�5���s�(� ŧR�˷�@@d<|/�S�J�͂�M���6��M�)u0�1�y�l:4i���Qm>�>s2�AU��#g��oy	���;��KH��^�Ss�T�{V�jQ�g$w��!7J��`�S�;*�S����A\���
�dS:�-���nCgZ`��҅�#��iQ�o�O���)֖-v��>�7�x����!6�=VH��~�I̡BkA"���55�������Yp'*�����OLX�.3jܹ�pV�4��/�n[�Hϫzk�>G&�ǳ>62{�ۻH,����n�2�Sx�\��������i?�<�EG@ �"dS:�K��� D#�� ��ɶC��Z�ֹp#"��Z
6��cnMZٗ�g`�,fӹ9o{G���2"c���`�4w���Ã�|y"U���ogt)WB��bS ��5If�
��r|ӎ�!FƸf���6ֆ.a7D\�I�[��p5j�	w��#6�g$�`֚���g�k��O�0k�ѳi�#Gߨ.]�u_)�4�)��u��>��09l}UbP#��S!��9���FkZA-��� ��Ϸ���Gh�LPGXʶ9�.��J����;����Yz������H��^'��i�pJi4��O�QZ|��d�����d�u��x<��6�W*�u`;[�C:ܛ%]��CC�|�Ix��眳�`��p���$���pߺu題^S������Ps���}"�M��H1Ӭ@�A^o�C^Ap��͏6���C�Y�
p�a՜0��/�;��!����^���ø�`�S�qJ+�t��������х�J�/�W�Q�VZ�_w���En���w�΍$��õ6<l�3����_4�d�s�[j��7�~9q�%�zB�l��d���A7������"'��}98Jd~B����i�OX['���"�Ы~R�د��� k;/��3+�h��e�#�$*s����.�0U )�&EPC���ӥ��zp[��{��"��l��y����w���=H���z�S�X!Ɍ�r�+H��Ԉ�a��^��]�������,X��=�>H�b��]Ժ�>ywf���EVe�.Z6폂^���S���s����C�{+�R|}B�.F	��$@M�|_[U��')6d�{bk ����\�����U/����
����q��s��;y���L� ��URu��|�'�6,&J�(/�z��0��a�eG���%
��J#�<ز�]�jK/':�4�c�r���(��	|��ߞ<����<�{�4[��4�������@�	˩Nw��ۼ�Z�����i��C���^�{���Z�v�_��	h��*���hU��5^#��c��$��������x���1��m(oJe\*+�E~�/{r�*>���)Ȏ9C���q�J���Y�q\�*s��\N����n���`���vت��(ɖ�q)�2:����6�I�f	6Vg��&�� �_#q�Y����CL�|�:��KΔ�Lz�%��q�
I؀0/@p�X��Z��˶K����s�*�IE\��]%���f���X�2}��l����It�ܲ8�O�1K%}:��$����B
1��x(�_�?�h�i�~�� u�c����b-���	FsMd�QI'��q�F�C����0űգc��D�}A��f��I���٭�l��K8R*'�Gȴ ��fP�K`��x�ۘ��(*�hjEac����8r����ī���_��3&���cT�9�R:�Ʊ��|����-�:SR��_�/�^��g�轠��/��,ƈ���uVtfZ��og#�zl�ӹ\8��YA�I3?�t8�lJ���W�o�Χ��/�K�A#3g���E��ʒ��1O/7�!�3P���a�"P^��(�(�k9ɧ@o�̂� ��mp3,��	��,6&G(ZVM������w�/kKc.��ge�ioW�������ϯ��P��ނ/��"{۔�3����urp��ϬW��I�Y!�U`J*n�љ	j�0E�/��.��nZ��MT�6�;�\�é�j� ܺ{����O.ナ��L6�[�q)�H�}�g_U��B�1\�}��rgo/NիCڔ���]Ze���m����n�j�9"�4�'uJ�R@o˒�_]�"��z/���.��Y7�Hj�ʽ��:�^O�5�`������D��8e�W7��c<p�ډ�X�ȪG?c��(jD�����&�;˵��������5^2V#����e>b����Sv�V@�J�v���C�-{�IQ���W���Q묪�pM]c=W-������g�[�1�Զ�w����&��.yR�2u3��#��̊nd��鬖t�BF� yk%R�Q�����dV�����䲊�\l�oB����6�d0{myF�:�f��n��QG�\>�i��o�:�	g]Cy#0о���K��f�8�S���TP3~���Aw�ۅ�7�V`f��Z�S��؛�&�rd�d-ǌ-��n��~`d]|��f �k�Q$�����c���-��'��=��سN4U���Xn���dܓ�̻5�k���D]5���lPgVY
o阻$��i������ɹ{���N�K��\9n�;υ��XW�&x�r�ش�2U$��6Փ���n!nSR�À����ns��}jiT��_NI@Zwk����%}'�H��O���c)��߲|Z95ٹʰu"]��XH�}�~Z3�Tg�%�f���o���%%�"�@����4����|�f�e@o2�lt�o��M�� l$QI'�K
�9�|m��! :������ L�7-�I�G*�ʤkxd�����#P��$7���4/���r���8B0t_эQV#a�K����u�:�4�n;��f>r�t0Ӻ2U<r��"��!��@��k4����=��=V��QD���P�f';X$q�������քb;�(�R������l5�ig�){h��S�Tǟr���_�4��v!��U�>��t�&f��/��A���jޞ3�٠}��:>���#���P� UoSo���%9r��ҷ2'��d��f;Ceu΀������-�E�*|+�gp�&��re�H�*��>78�6��?�*�������W�����r��L��m.��?�	D��7�$���f��O���L,���n�2���0��D
�:[��^����OjJI��Ҙ#�������#6��ƿ�my. d�ӡ��U�&<x5Z�E@Ǫ��y���v� �F%E��EZt�]wuZW��;%T�����/�P��ʟ��Y�(q�Z�l��_ql�ycE�H�!3/�:����������|�8�>���BҮ<�3 �Y�c�F��H%���CE�o�J_��t�a��S���&g�[<r(\�?cM��!� Ά�?�4h;�?	��G[�f�$<���lg��5���vy�Sh�O��v�~iY�m�L��:*5�
����6��_��{�b������@Y'&�y�F�vs�����6=�)���+�a�����|�����K�p��㴮�k���zv.s���5���h�.t䕻U�:s���ͪİ�v���[4s� z���/Ђ� q��(�ƘqH��G	ԏ���r�[4���6m�rb(�`����*.�֏���bǔ�oTonc��w��}*V���<Lj�9r"���F��2+w1��|c!U�.t�n�#Qj�s�l�v�)�T���O~މn�?��RQɨі��#%$��/}C+_I�,'Һ�%�@��J���f]�8:tm�cX$+��ڰ �.}r��<(��k�CF���8��]�Ҡ�AL�)� �A�sV��>2���Qז�R��d$�&�`�Dt�QQ(�u��eҭ��V$��&:H��h��Q���>ՐUJ!4� g�~@y��{�O9�K��Z�r�!S*T�DsxV�{��U� 7^ו``�&OrSH3��U���lJ�dgl�-��nWnY`^���-�9e�Q�଺�"�=�-
۲�R���� �(I�Q�v��|um�56�kU�->"�5�Ɗc���Yc	��������B����V��.��E��C��n�a$Ͽ����&2�}��o 2�>���6⼪i1n�S�6ŀr.2�(���w~iSJ�ى�@"���J�_�����	 �]���Z�J���u�"WL�4��.�Z�j�g��8f��o7�� "��K��2�4����*\|������o�U�t=h��G�H �3�I���
���|gl�!ZV!�G�����7X�)Ix�����r;~#�gE$���.�}��4����c2;0��w�ǡt#�Q4�B�u�XZ4�K�	�Z>,��0�EUv\"4!�,�:s�kn7<�T�������K)��+'l��2�X�뵊�ޞ�s�P��;�;��Lۆ̡j�eR��#�,)���h�Z]����r�p���;�ng�v�{�Up�+>�Wz�`�ͱ����F�x���V�S:2���>���#��P��Mo����"j9�޶�L+���{�^T����@e�n-���㘬X��B�*�Yǉ!m(�7�.��e"�7*r�(79�6�/\?"R��L�����TW���,��L�Obmh��?��uDz$�5n�V��l~��Ѩ�L&:���ێެ�0��j����Y���^y-h� 4j�7*�LNG��t9�����]���j�U�'�� ^6l� _��-��x���E:�阼�D�%��� �pM%���7��ZQ9>;_��_C�\�J��\ǧ��(+��Z�v�ר�l+���*��@�tJ^�(S�@r����!8W�Ӂy\#B�H��-ѫY�SF.��%]�=Po��X�7��u<S�>��`�.[�C�\dT	{�-9J H�W?��h5T	���[���m?���S�l���5
Ӓv3��h�.Ӎ+c1���#Y~����-5�	���9�X7�K���w�y�|��fD'`����N�sA�����=��2aw�{a�I���T�������~�]��Ko����{7fv(M�Ou�m�J..4��O�d:��vÏ�$�ji�v�}[n&��§�A{�|��q����@`�H\ŚA����Sb�?������1L�G��b�{��Tį*(u~wU�*�/b�2"o	�.n��yw����7�*PD�X+l<Ƽ���)%��������w�S>|&�(����Q�D7Q>(��[) �����	��ރd�?�Q/QCE��
�#�e�i?�+�R�,�
=��	��=�R	��841�ٝ�@+r����
�}l��<bj����Fh�h8��]�Ȋʻ	�)�a�;�Ys�3���ʻאN����߇�j`f�ʒK�O���=�;��C0��Y�:��ߔwI�3�p1�Op�)��A��z[������do~RC]�uFO���p��������0�^�	
�����ҔǛ0FӋo+?cYX��Kw��?�[�A����P���v���j|�m�/�*�ՠ�������2E9A�Q6���&{ۀ[�m�B2f��?���>���G����2��G�_���!5�����T��[u�G��L���_5&ظ�b!����Q�T� ���擿��v����{N�I&!>�f~r�e�r2�
��g<��Ѯ��4�����s�;���8��6��$�)��SXM�(�)���8]yR�-=�h�>�N�wƙb���C���"�������ѦJ,j��ۅ0�Ib�����tv�B}�H���B�{���#����#�u@�,��L�AJ�V��⥾a=��NE��-UJy6�xw�~��c����ZF[-���>6IcU$Fd������M�(+.hG���p��2+�c����u�
���#t�=u��~�=�pu5�s���0af��Ni��m�= �4X���M7,�����݀P/��X�;S>{�~$�&E��kpGviVP��/%��F����$�]N��k�f&��m]~QH��c����6�üخB����^���+�~��c@���� �G�q�y���˗j�P��z���#�Q���b�z��g3��e� j����V2�}�{�MjTw��vC��?� ���2�a����1DqP6��2v�7��=r�U��e���I[�]:Y7\�v댡ʅ1�{7���a���®G\{�Y�]���z�+�����&y3�!t4�� � iC� ���Ћ��{@Y���c��3� ��"}��G!D����N���@7��e";���Ů1�S��,�}{��C���oWx��kI�����Yh�ܡ����ZE��KR��־�����@��3��9a�xW ��`���(���J�e����e�RN��ǯĂ��sR%��Ǔ+���������WRN���3qc�`�������II��B���� !_��i��$rTu�ܸ���ܨv`��N�:�|Ǚq�,�5���N�u8��:J��G�1�F�C�O��Ь~.`�)gc�[,G���\�I�}���O=͂T��ԡ�55�
�Q)�c_��4T\ E/F��j2v�.T��C ��e;)Y��n��=�
/�z���Q^���7Ȏ�1,`���+�?�x���\_����`�Uܘ@͈�ݪ���:�&e5�P�������j��KS��������<������2M�Ѩ�8�jk���~�|���Gk=�e��� ��6�(�_4	�g�Hk,ɑ��R�>ić��i�@GVLw�5=57�����Cփ
�cZ�����k�ȆlTBh��b�0�wO*G�x�R��ak�,��m!K��uu|���E�}�����xE�ŝ�hr
G��i�K�Җ㰳S��E㔷
O���~�u$�S�Z��`����7Ĥk�c����,Up�M��j�J�$��q�8�;H���u��n��,_��G���Z����js�=q�sh�>��I�yJJ�p���Ժ�Q�.�k ���F������V'0�o=���X�A�%����mh �e�����_�Լ{t��rPi(��g�:���Ķǭ`�ry/#EO~ٹ��D;��:�n���tL����e7��K��)L�y{���Gcٺc�|�Ta:��"i�ᔦmF9|&_�b�+�%�cO�r�a�Bd����3I�I��S�;���<��}�ѳf��5 ��Oa�Hn�G�<F;p69�zaX�.�*Lfq�kĻV��<H���m`ӵ��e69k�x��m���&N�*�x���v歒���pF@Ӣ-�f�"7���S~6���,�����%�#��A�m��,^��m�Ӊ��];� 玐��mU�VQ��^�N��+'����b���<��5�V�g�;��hV���9ΰ��kQ��q�(� .�)\��ε9}��F�Ү!�C �ռe�B�C���L
���M}��(B@OB2N�NcWwS��D
�~o��'E+�p�	dò�hW|�\
n㩱U�L�w1%J�q�d�N	5L
�1����ξ씃g��1d��v�r����^tj&��P(�h�]��c�S��3��e�r�G�c�G�]�.��A�ŰR&e&�#j=�'���	�rD 
S��V�x�R����	����� ����@�r4Kq������#ӝ��r~��T��V�`��պ�P�����KpZ� ����q�� ^C=�>&���߶Ι�	����kwN���$scQ�t���&\�r��8�S�WN��T��!�7Usħ'�U��p�z��pJM�n�g�M�r�/��d#�#Vq�r���t��vM����~�Au~���'jQ��������P?޽a��_��t�4�/�U�~�'?�W,'�Iyh=J�ݾ���²7�4$��٭���Ģ��Ϛ�s����1��F�bq�f�cR��U��]��Jt���t�s�i}�����n�+pC��ҹ��`�Z-��<�'N��B�����1�rzfC�d�%B;��#��9�cۣzݤ��f҆_���J���B��
�fhTT�������!f�7�x�H崔]�I�k}M N�riM�*�UӜ��iA��.�A��L6�^�W X�iD�֮Ԙ�;�٢���sC���DQ�����o��d��'�$�Ps�z���C�	���1�w�2TЙ��^���PaH7u���	�A;���d���	��h⧒q��j�c�!�,x����@�_�e����[���!��%$c3��>��t+I�`�.K��:�ؒw�������;up�#^��n��W��dW�����x"��	����U�^օ�C��Np�x�=bm�*��Yd2��c0!�����hg�z��/�� �=���JҮ���]5�3����i�J���W�
�V�/�_Q�����gw�/P$Oül��r����_�y�d!�µ�~B�9����(�lگ#+���3��n�5ƅY�'!�O9_Bx~I�x�z\�ܩa�m��Ɖ
�Ÿ������ǩ Rи�x7���m��e>�$q0F��d�.�[7 MNEL�[��8uTzuB�[���&S��D��~�~��`�Ǐ�6Hk�z��ߟ����F&+O�d�oj��L0�6^̠S�X?���eS�b��ԡ3jy��f*ǏE݀�.�¤��wE���Gs�c��x��{��1|�u.�`V�Y@t`_b�׈酬)��E{�% .K��I׏�� UVX����7ୃ��U}�y^���h�1�g�oUy\��HZ'�i&�/q��y����.�G�d[�L(��Q�<���]�+�/��4��ҁ�c��o�8	�G%���<�,��%s��띭�;іl����c�	:W*N~�mۣ1�Z�:C�k����;��@,�{V�b���:��a����<Ih܅a5�gX��4۽K�����~�)`4_�������J��+8n��V��1�y��@r��,0�����J����X�\�����j�~(��5�����p���(m�qP52A<H��;{I��6�A
V���=�_jK�q�/&����C3�;� "Ku&8LRE�C	�Ǝt���/G"�Xh�.�U	K.�W���O��%\*�P%��<f���X��!}��Y��^I�خ��`�xOl%��!�+�P��/�	���/wL���.T��y� 4��F <�^O���h��Ͱ�r��}�]ޱ:S���7F�Y�8r�JE<ô~2���Q�":�a�����L���k��򲵂����z�F���s�MUa33�"�� ��=k9�V�&�W�C'���5xO�N�a�����*(3���.t�;@ �<*�0l��/� �S�h�H�ӏ�r��;����d��M�L?ߚd��V��rHG�m����Bc59�W���!�}�bG��,ɦ�#F��~�u&p�u�����"Ŵڠ/S�����ɡ?^��;�z����A��`�����Q����x��¡y���	�m���V
Wo�7�b�G��Dy�!Ȥ����Y���p�V�K.;l�hOй���i�.�uQ�+3���(Bz@������H}�4:��,��|A���B,�:�q
�����lK}�}�B7�lO{��NK �W�/d�݊�
�]oo�pS ����N�d�ET�kb�W�&�\�bZ�j�l�%_~1j ��
6d��"	��v����oqY���]@�1]6%v_�1f�� Y�=O'W?�!�U�\t�L&Y�L��&tB��U�\����]N������Ŭ&~�M\�4=�)�����	��r�KS�(�q����<ٷB�ƶ���1�p@L��r�XמzT����#�c^̫�Z*�������8�P�u���Z���Uidq��^�9�=�E+&�!j������¸�8|�k�)��#4s��6tM&x����8���Wg�f���! ïs=�����?�)G��� =M@����#��å9O�iq����޻�ϩM�>�q�zˣ$�'�˨*�6ژ�8?��B���d��pz4ˮ�U�|'��D,�2�y!�I��������<�4]M�V��==p�\��,{������F�p�ӟ��R ��Ea��懎x:�s�毠��r��D�dj���!ێo`mVH-uJ�m���C���-�j�˛vz�;����B��#_��\�`z��q�!�q������y�B�Lw�?@YT�nG� ��Z�㽐�g�������q�$�g '��iF�*�����&�Ak^!./R{l��"7W��#i=xǮ�ܮ;��P�L��CeD�ex�K����@��
'�q�P�մ��WCPb��[	��0[�T���qv^��LP�au����1U�A��_���/�o`6z�-�����8P�+g���"x7Y��?�:8<����[��Z-G%}55�:\��@�I�z����3	i�������?����u	�N^s��1���p`��Δ�"	/�h��`4�^�7�C~��p�|��V��c�Y��~��N�0�{H�[�AW��g�'�%�9��s�JKpU�Ny�7y��?�J�|�W�B�V1o�_�{��eK�;/jw�s�$}�գ�l�D���:�_$#d�}�{��WO�9�`\����l:6����a0w���>X'��~9XӁ~b��.�5�I"qXG�n�B�x��W���q8�0�� ��"�њ�#l���M�e�$$J�/����.� IR�Ep����,�ћ�z.<�[���r���\��*��V��?`H}pz����x���{�+h��Ԩ���Sc�}?��9��9XH��^qMb��ڳ�y8�}f�9�EvB.z�0��P��{��-�s����x5{K��|�?.f��/T;@m l_{�a�"Xt)V�{4[* �n���²qUO1~��L��2�����*qy�X�!�m�@�)Ur��I)'�&j��/���(��eG��Eӿ�j0<�C]�/G�h40Ys�����H,�	��j����<���\b��T��T3_�%�����	3�\N�����ЬZ�����+�c�����6{/�zȰ�5�?�)Y�J�~㵻�hu�55~����ؽDD���)�����L�7
4�%+J��e+.�O��J�o��Z/�.���;zx��J�g��y��\���	Ϥ�k�Ŏ?\���������e(雙qI?�2Z�����I���6v�����@3_CC�q�"����Cl��Z<jK��L�����z�O��i5/`}XX�O>���K�-PГ?N�iX�\:�%��Zf��X��}�Y�kXI��۲X�%�Q��%�c��D4r�=�~�b���1ˀ�9����#z�@��c�Z��س-�R7�)Mma�Qi�ې�6��f<��$&U�a%���ɞ>�}a�,f�e��;|R��z��1u�k��*G���gp�@�{fp�K��x����n���#a����Q�8"�������滍��S���������RZ�
m��4��%C�Z<�R�$3_��]^ԏg.{`��=x�p�:�,���t�+��7�tgC�?l��*�|�L�y�UA�r�_.�tXq�j��	M3����:A/��pAC|���a۽��M"Q(BW���S��xC�B�x��(����Ǖ���� �}m���,�n�ĵ6F�y(&��M�l��1 �'|�OL�c"3�����<u����L����vP�^�OK�B�����@3Ԃ�ܕ��3ӟ�̰��i't! ;�`jo��j	>��Ov�N�snzm�M.��63=ŗ|@u�(�H�@	Z{�Wa�o#�����	�6��h��xH�Tg]_��3!J`gfek�F�h'��-d�"�-2��nZ�@`�c���8	�\}�Qa�;��ϑ��%�-�L��U?�oP���2�ѳ��Ԋ�~\,YI��ؚkX���;�5���J��Y�u��8��C�E��xaʦ�܅�h�nҧ�����uV�&5���5�n2R�»��-ҹn��S��	�l	�+ì��Ni�����i@�]��60̢欕7��e$��}��ܒdZ�����":+\a�镚RSZ��gW�<f�FCo2B��b��"�[�!��4��
���|p��bBZo��t���*�0 ��ID��
�=>|�j1!!Wk�$����-7�J�IҎ���u��[�#���$t����O��袍Kf30b	lъ��#�ZӨ�7u�6�4�\����>/��00]9U9`]¿��!7���k�d	��qa���Ϯ�O��=��""Xa�n��"r�YԮ��O;���XO��B׈��ܦ��)�Qh	��q�r�����(Q�1�nv�P	U�<�>�������0=��I@M��o��@��v�]�*.>�j#@�P��Voq��Y�!9oAa�o�dJ�AdR���e���������A�*�L��_S�pz��q%Me�J*u �7v5e6���?E��ϸu��IXW�Y�i\�/s_L_�#m+H�?��`D��q��nЙr�����JL���񵊻���1�ɦ���t;�n�^|�{�c�jG���oH��P�5���������*s� ��R��3��P#Mxr��E_�,��"���� _�%B������Z4�Q;�я�}��_z]���Ҟ�V���UG(�q:Z���M0l� �x�~�g�7Xa�Kַ��������8�^�|�B�\���eCY�t�FQ0}%�� �o����IY��zSS���#%�[���\�G��X�p�h �A?���h�y�	�	�[�����B�h��l�F5���v6��h�΍���YyF�g��B	l5����&U��\�ꉐ���§@�'��l�c-�sD�d��=���U���a�V}�
����3����$�`�Bj&���iv�p�\���n.1��Ye:pd�ò)��Tv��[��9�8�>������Bq�b��c1\Hߺ�$=���u����^�Ma�
�{bſ��׌�*N�Sl<��m�b���ol;�n`}�w�OU���*3P'���	<iM���E��ե���w�}�|��"�O;�Q��QT6���w%)����U-���M�f��?% �Q�{n��U6#�2Ǣ,W#+�bd,d���H�a@Q��r?��8����`��+�B�=�}O`�<�>�9�FkǄ8�+I]�g���)�C���sӚ[l�ʾT �����Eiߪ&h`�Xu�.�K������C���|Э�<p߷S��'1�D�p;�/����z^���F��'��~u��]��F2��]���+����w���8
Y�ē�n.�J�F�b�+�IX#2w�頾j�Au�6�������5���em�>��-o����=œ��2h᪑��|��c���4�mXD�2i,W?��>���GAȇOk��� _��)׫�62T\2Ou��=G�$L=j��B������!�z���-T`��۾0�����\�mQ���!��af���pt�r��t���������ٿ�|��@��>-�V�����G�
�JVM�.�&�[�"M�`N�|��- `�a*��d�b�*�C$�0�ŕw���b�RB~�a����0�%�buO��$�.t&���B���p�,���#=�3����@,�J��tJ�$�E4�a �Nh�&-�al��w���^���{/[�����cxJ�dg��m:e��(έgG�;�p]��i5c���Tʵq�t=�=~[pk�����a������*\=� r�*����O���{���Tu/�I�ޫ�{ �R$k��E�Х^��}�i9W�����^�C9$��ɔ8)��q�&wZ~4�ߦ%x�Q�6��L�B~��ˁZW̝K~pr�c���K�G�#R��ԼyR��˺�~P�M]3��fs�}��3�����(�j��	ɗ7�2�P�5ǀ��$�j bwqGlv
kq� ��2|gB���D[D��E���ͭ�h���m�p�%�܂�ݲ�Y�4�(��/1��4�����.G�c/Y�NG��)+��jx�3���4D�l��)�caB�8�T�a@�-Y�&B�3�����D/%6S��N�x�@�e�J��5g1�Ú�{�Ny����rU��(*�ުC��A߅ha$J��'���y���ӬKU��907[�%�֖��n9��x]^�G��"v�|�@�h9e@�N�h:�ݏ����􍓎�ǿߛ�ޭ�ZrNǚ�3�P�`��<�D�ԜIk�?��a ���m�g�u�e	��u>�ٝ8��D:�����GK�l��b�u�:M�GP"PF�@�O�~��/� C5Cg�:�ϵ��D\I�z}W��O`�*Tm�}�s���M�o)E�D����\����h�ͱ3U�&���1)���n��z�m8�z��>���WN��D�t���c n�B��O~��P/#���U��0{��M���n�~s5��ۢ�hKWzj�f�K���x*P���M���ήC�����8nK�jN0���|T��J�������%�YU���]�	g67H�ד����R�Ƌ��0iF�+Vo�l5�w.(��Q�ֆ�Rc��u��(�ki�l���8\���0�O-u�xATD��k�?��𘨽j݁|(_3Esju��+x�D���6�
j4�i�C�y~����$E�t�
Rb����8/v��~��ɸ�7/S�I6����,�w,M���öh$*�wqʗ;�~e$��;��q
w,�σ�
%���쀝>Y�M�u���2�!�>��8�|�J|���@ m�=e���kEc��N�(����G5�؛����X?��%�9K�>(�;� ���7��7��rs���G�Y:}Sd ���r|��f��~�&�gƽ;�~:�n��_��L�)��~���ǵ�������0*�ٝ�S�><a�<�"l5�	Z\9?��&�&�-˿�W�O	��aL� �۳3�U���ߋ;���<s��L�U@a lqORs�H����� ;��G���5���L����V��H7 m#����O�9�!/�����"�4��0��MY��pW���k�p�A���X(�o���'S�A��旗��������A�҅�o�ɚ�L������Y������Wm���V4�!���`���.�w�K�5%�`��O�Z�VV�2X;��Vh�)���=��X3QQ���>�(,n-�Z��pB}��f��B��7���mB�����
Ե��7�}N�fB!�<O��N��2W�bY���
��{o`���-ʻs��d&P�ձ�W�cg\�4L����S,1����2d�n�	��|�T���Y�K��^���1�%v�_�[�h�!������۾K�~���Q���W�6�P=�5��4��^�]x^����he&ho����=L���/�N	��r'��S�D��[ê�'�l�жi7]��J�@6,r���ā�#֌i��Mq�qe��Ȋ;��@���P ���e�	Z�bM�9%q|��^f�#=�&��
�"/r�����"9Mkڃ��Ӏs�kqt79�&?׹'�8d�VWQ�����,!�,�s�4}��.�S0h�2�M�<�j�ǀ�t�l�#�q�w��ꍋ�(�MY$��������'�Đ����?!�}���U�4�0�U~��'b��,�|�yK8<� 9s 2µkz4�Y��p�V�����FM��Vo�
[���F����HbRj6!��)���뎢Տs�悠A쥿�H�莊؉N9��8�d`W~�-�o���7��[/��(#蔻�5�#z2[���3Bv�#ɖ���z�$s�K睆"�Џ�o�c�1Bޅ����>T:����a���n��&J�k}�����N� ���i� 4*�{���nwAի].�L�e�x�AofWc�<i�����;)sV����C�i�D����uqG�7�-�ʳ'��P�1����C�p��E��Z��x�N���k�D�!�����B��@�3�b
��,�X@�ϑ�$��q�!�)`�٩6��j�2���%�s_�n?tPM���68	E�!��m���%Y{?�A��:�o�(�B~G6��b6вHU��gd|��,/�1�q\�������ڔQ)�]�y����ZW�����"�́���wL3�W8�]j�w"�dg/9".�=�7�2�O~�_OkO`�����F����D�+e��7�۟<�������o�&�6��h�D<�<��D�� ���\6���iV�ÚyV(P��{b��:�8"i�8ƕ�oz�fﲰ���N)-�cy�������pҁ^=|���i����`���yvc��ʊ� ��r�R=�3X;��wy�s)��@~ ����'� ��R۰��H)Td�x��d��g͡
S���ߤ����[I�0@IVy���:�䰬��Q�>r� h	_�g";�y����D�KN�c�}�YSrRcT����(����@x7���`كZWS��� Mͥ�=d��U-z��n���`	��8�i�&kQ��E��՛ȩ�-�Y<�����τ���%��%˺�?[���� p�k�H���5�<��Q��eY/!阀��α���H[[���Y�3����n��J��ύ�&}�+�}�c2�jR��u�u�:nFʾSp��]�d�s�m�"��i^ݻDr�@��#:���R���W�T[����$�Zn��OB"��X�#����Z8i�g���f�^�ozc�/�""��i}>4�P��"D�|��2��"�o��t/��r6� 1هI�%Y
�3�|*x!e�ue��l}�EQ�7��FIc*M����t�&��#5w�$����Y�������j���0�X���ʫ#F�P��\u�4S���r>w.�0xtDU�`����!fL&�e��k�H��?߂�B$���ҁ�62�K�HX��o��e�ל;��;�������[���M/��d)&)hQ"�����r�F��9���y��v��U;ǥ>��4���ױx������,�#a�����r��>��#��P��oX�s����9�)���׎�+b݉�m�+��e�X�	ї�Wi��M�b*aA���A��cӹ��eh#*�ƈ7��g6�0�?�tr�c��(=!WJ?A�N/�w�L�VEms��?�5DE*ϑI�z��CW���!(LѻW���G� �yy��Eqd`���^��N���j���!2���~��߀��6��U:�rY� 	���̞�ģx��Eerqt��/(��k �c%�5�*z��1Z|�8;�R�JJ�������+ƞ�>�(�� Z��E�bY�l��J�ƒ)�Hd����+��&U8��o�d�@B�bd��4Y�,�F���%(�hDPoL.a��n��f��S���k��[!yX\/�o4����� 3x�?�RTh�ش	�QX[���8�F����l,��5��8v~�Phf��6��c�tYI�}¯J   ^   Ĵ���	��Z �vi��:'��(3��H��R�
O�ظ2a$?�K&����4`��̏;Y�����,�P���#j��6��¦�޴J�������'��Ɲ����dL�KOZ��P*~�n��ѥ[�$K8O����7;�b�O�I� [�8IH����5�D5��I�=^�;�M�LyR��	�Ay���0��	D�+�t�т�/���`옅a��W�o*X��p$�j���Ċ�<j���^}b��"e��2d+!�ĕ(ǂ�1mȮ&�"��xrd0hK�yZD��tf@8=���2�'�9c��9E�8tp��с\
��O��"�(O���N>��&�8� t�d]��P�D��<��=��"<1�AD-0l��u�$FgN�i���j]�`���4L��I�V� ��P�W�\%��Ɓ"hi��'QjEEx�/�R��� ������=&�ć��1m�%��(�t��3%h�A���4��b��Ƞ@O�U��%5�	�bj������D��R$kx���ʲN��a�j�<i��5C-�㟰l�]���#�>�F�8wA�p>�t���	�n��,�|T�$XG��/$�4���'���DxrKc�I4/�t²*I?��\Q��*2r�ɩU���9E�Ʉ ��Y��"P��˦&B)nN2�Ę%n.���NS��3�a(�]�Jis0�.а���	n���E�L!^�l�+#Q���&o�0�H�Od�����?��'��D���L�(=f����t�8�g0��,zJ>yw�\���T�<��퇱 B��D� &@ܼ��%K�7�P��'�ղ@ ��G�!�$k� �  �                                                                                                                                                                                                                                                                                                                                                                                                                                      C  4  �  ?  �"  �(  *   Ĵ���	����Z�/C�'ll\�0�|r�'a�	�Dط8��0b�
�<�}#�'�t4��B�h�d�w,�:?������i"x�	�-��K����1Bʚ�HH�� Ҕz�J�[�.�0�|)`��u�(��dů,�HP9Q��#,��5˃ݕF4�,��	�a�l"�i_�6��	�aι ��0xЅ�)8���ڛZp2�"n�}����D�
�ZZ�Q�W��".ٲ�0V��	DWC[*~��?ѧ�ϔ&��g�WK��ؑ7�Lw؟��G�i��)p�ىH'N�1�Kò
�qK����B��B��};�6	Veg8D������O^��Eό�	0
)9O~���<���H"��^ӔA���QN�<	��A�<�>��t�)��"V˟F}�a݄cx0�J5�%��S�*h"`�5jO�2��	�uD	�w7B�bajE[G�Ď@�����L�8	�OLc���*m�]��ɤ!\��*ыUu��y�N�?O�:���K�	�B���гJ��4��~�0��Ǆ�B�	Qa��p�I�0��рg�
�"?	씛b����#�8'���ҫ̸X<�9o��yB�J�x��c��e�,���ܣ���H_�-�{���2�|M���T�x7��Za��1P!�$�3#���7��$��I ���%J�'�\\�f�Ix�p�Qǘ�$϶�@�O�ک�ҧ9�O�5ᄫ�1�����Ƅ�m�LS �ڵ&#Ш�ȓC@���VƇ�78JUQ�O�A��D~2%W�O϶�@o��*��ң���B�'ArA��^� yJWj�$D�^���'rf<r��O�Z�iw�C�@m���'�x�+�%S�t�G$�N�2�'��h��f&��ݥY�paS(2D�xI$k�X���yA �0j�lK�)5D�T$�K�m��0��28�딀���y��� �X�3sl޻b��D5�y��z�S��.n��isjO �y��B�m[rCU���\�KΟ�y�ɘ�����Џ�p�����Py�'��.��怛�)c�"�]�<1������q��I�:���QY�<�0���(�~ 8b[7e�m��,�X�<���vR:DY���fɖI�P��x�<Q���1��i�edH@�,]J�<10C�$b�89S �n�B���%
%D�ܹ�l*5d�x�w��l�pe��>D��#p�����- v����0D��k�U��T�����|mc��?D�0Ӧ'�9�
����B��(>D�|�$@ثg��@�E�*l ɛ&B)D�r1MF�s�ᴌ³ �<#%�6D�t�I�%&ԉ�gՖ��$��M4D��1S#� 7)���';��ՃVa0D�faR(:�4^�L�����B�	�2���@L"_��`��ڥ[��B� �|��	,p��PEÙ=�B�	4)�֩Z��8X��i#H�9��B�	h�OV?"x* ɐf�`ʢC䉛	�89�bC��00�@A)vB�*O�,i�,G��ԳQÀ�DJB�I[����g�4Y��C�K��! 2B� /��䉷L�57���sD�$L�B�ʢl�s� I�Ti �۫*FC�I;@��L���2?䜀 C��4�*C�	�[�:*�ȏ7+�xe�! �\�C�I�`@��iɄ$�T��s��%�0C�	�p>\&��%k�,��q,K�O�C䉋
̙iUg��t���j���C�	(>�ꭙ��U�u��QJ���,�C�I[�jh���:��	�V(�'j<8B�)� �DHG9&P�� �� =��"O��SQ�����c �	�"OB�c�gG�[�~h
 �Dh8�#"O`�A�L6��gfl��+w"O�9�ΐ}r�/��|#�n_2Vu!��L%~�.A�UHU�^Q�"��+kT!�d@���Ekg�B��Hrb�^�DR!�d�*�~����H��$Rc%�0(!�ā-[�d]Z0���9zAq���(L<!�N���@���%%D���`�P!!��8�@	�Ī�n�Ij��{2!�D_ +���A��4k>Kq"ؐ&!�D��y0P��M1eH,����N�p�!��2kr��z���dA�����:�!��/wSx��M�Z����5��	Q8!���}�p��#)_]�T�P�RM+!�٘fi~��.�.���i��V
KC!��b�
�Y ��B�nX3$��$.�!�ėua��0��#���*��"m!�D�5��X;7�1:�12��(?�!��`tȸ�v אN%�T
1�e�!�d 2����HڟY�e�'l�3~P!�$�!-�ԨhV���i఻�`ɿ"�!�Dr0};r�۷V"4[ �Y�E!��U�:�J�# �UAD�2�!�A6���&�.aը��k���!��NP8X!��[rĘ��F���!򤁃fr��ڇ�N#/O�|�Hާs2!��T�,��nO��cT��9V@!��,@n�5��훌#�֠8�M}�!�Ę�+D=��	Y�Q��Ղ�JՓ.+!�N�A4JA���P�W�b1�ႋ?.�!��9Q숈������L�D�!�DC�p��tIO�OL`�3��,3�!�>X �P�v��> ��r�@'l}!�+n�h��%Lz��Ձ3��y�!��-`{J��� C?N�\ݲ��7'�!�$*.�Xy��� �/��TS3��h�!�DQ�!��y�"�8�8I e׫e�!���.�E�ǟn�MrS�Zi�!򤔝=|1���+�IP�
]u�!�$@/̎�(m64�K�
7�!�pM���Q��X�T���7�!�DM�^�\=��䖃u偐�Ƥ0�!�Նin"i3��X��R��6�!�:�J��W��?}�}P�Y�:�!�D�%ei�|�1�	nϼ�rS�A2�!��<�4�٣�	LǌY�d �9!�!��7*��g��T��1��:?H!�$�X��
ƌƭ3������%+�!�$���t��u�Pjw�a!�D�=��q�'OC)m"�,�ƅ��^a!��΍�v�jpe!'`p!N�~B��w�h{wg�)#� ��S.^�дˁ���W7�3pH	������%\O�<Q���x�pm�ѣ̳-�R(���%�E�6]��=�f)�i"6�ɽ~���3Ee,5�@�9�oْєB�I#+P���/UYv�HTR�V����<]��ȳ��P����㤁;�6�S�\�b�hEeã/�¤;%#<FwxB�I8.P$�:�m�t�4G�l��Mҍ�
am�c�n�⠎M�IKK�08��r� �,]A�CNժFZL���s�@�ђ�9���;�KU�m*�͚�	ۗ	�z��G��s8T�ڢ�׼�p=!7,[��2t�d	��[Պp��x�'�2%�T%S�	�H�Q�q��!۴$R��HJO`���fU�DE����'�^d�ea[�+XB$U���-y�'�j\�*و��y�e��2���t�π ����!CN�������\�a"O1�S���BHp�0�%۱�}�!�E"�4'�p0ǉJ�]�')qO"tcs���r��X�-[4F�|J��'��-�ԅݙgl����k�/�$)�δ%JԱy���o9V�0�[�R�j���O=|l��W E�Y/���d�R1g�Q�����Ν?�P%�����.q�_<��AIR^�(1��`���+6"O�U���n����A!:V� ��O0u��aT8G�
�#���z�H�EKW�O��z��͗ l(�����2�@-��'f�0hQ�Թ2H� Ɇc�z�X4�g��V5L�)���Lx�����U��	��'�(h9R�B�"ItR�K6(�j
�j�������r��,qCW�o�\ ̐�0�f�+��"Q�t���I�%@�z⁚
�<}ReC6NC�OX�O(ɠ��ۗ`�6e�u�4x��≊<
]Pp��J�?_D���,�kw�a�	�'�`�c�H�!�la2���g.a�'ڌi�e�	��9�ta#%0�H��8ʧ��xdO�BRJ�0[���H9x�h�)B�z\v9���U%�������f"ը�i��
��U���\���~ܓ��<3ҀѼ�V�p��\������	�C+��;�h�U�d�B@����Ue��W�6�R�GF�l� u;�_�p=�TGν=��T�a�ֆ<���
h�'5d��qNG\Fjl�7���:,`��ش{�m6jJ����3��R�f��`��'I������.�0I��D�. T��'w u�Mh�Rtk�Z�d_�@P�t�O�|d f�̬�n 2�Ǆrd��j
�'�dŚ6�84�L1{B���$M���BF�)�p�A!�i��s��١P��'s�qO�б�R�<�D�)R��3/:����'=�ěDD�
P�h�JV�U����OQ�<�|���F�$�l`RU�ԝ����$MNE���� ��\���ܟ�Q�`���\�KH^	��5L�H��".}�8\�W�#�4�RqH��X��U)>D�8�uc�X�kb�Qh� pj��>D��F��d����#aP6'�H�;D����	��D�HQ\�ę���'2-!���@���@UHF)}m0��Tɘ�,!�$�Q��`�
�}�|��Rm !�$�:3�e�1}ǌ\�RC�;8!�$��<��U��>N��i�B5$!��&*r�J�!P�����q�
qf!��5�ݛ"NԌ��A��T+!�D�1b_���� ��l���mG!�D#k���s@��XW0���B
z�!�d�0Ν;e���:U�-CV.�+N�!򤄥r<d������>N�L�⭚%�!���8j"<�`k�7'S���fAu:!�DT&2�ڐ���Ǽ�e�&c �z�!��܌d��+�!_�[���s�B�}�!��/O�-XΌ�~P����<(!���$h�zte��d)�H��J&n!��Y<"
A�E+�+$��wꗍk!��M�gs��x�Y�kd�C��4�!���<\� �$�ڃN�d�S�
���!�$��F��0/[\�"����!�D�T�Ѳ��L��-�s��Y�!�]�)<��@d&�E�U
�n�T9!��&.�8$JP�[�v� �!a��_�!򴴭��_�2C���ZD];�'��鸕hϷ]��i^L��3
�'2(��W�.����gͻG=شQ�'�`��%6�2���͆�&�'�b��(Q+�R�6���dԕ�y-IbRj�ڑ/^%���μ�y�,^>_�<�b�p] Xh�+�y2J�3�KƱj��KbCC�&%����RTr���C�Ub��
x��	�ȓ ��Q�ӤIrT����1_�(��ȓ���ٵm��
!:� �#~�&<��t��舒,J�x���C�ܿQ�Dن�S�? �{u�۠���kA�LJ�sC"O@%#���%:p�9r�AހX��9��"O`xZç�=��*�*��@����"O�`�6�XM���p3���"O\�E �N���d"L-N8=:1"O�8��g�!�r��w��Jl̀a�"OZĺq��	Q7v�q&�N�iǼ���"O�8�uĊ$a��H�-T�/�|��"O� @R��$o���gÌ$f���( �UH�l	xX�h���S$S��ɧ�Ũ��՚��,D�\���!0����b*1>l�zF?D�����ljj��em]�,uHi�7�<D��Zqͩ0�Z+]3P�}���:D�s�łc�j��'<�褰Gk7D�\BFE�U! �S*D�k�<1+D�h�#*@-Dڼ% &GE<�r�)D�l�WN�(V>0b�GV�EP��Y �;D�x��-��|�蠊j������:D�(�F(�U��(1��+ *.]0*:D��y%FZ�|XQ#�Jc��c!�7D��(WMS� ���Q.
�-�����!7D�P�$GC�5j��
a5~�Bi!D�ha�7o89wa��vNNm3�:D��A%.��E>q�֡F�~\!b��8D��e�R#wl�C2LÈXi"�Q� 6D�tC �� I<1ڇa��0A�P�'�8D���rM=I����T��R�(6D�@�iҢ��eJ��3/���3D��#��՟Ql$�[��[�P��	?D�HBu%^�[}h=��9?ޥ��@<D�����J<# ���o��후 ;D��C��+^m��C
,yx1`�O6D��hW	U �P���{DC2�'D��vA�>� 8t�����!��#D��Z�ꎱ���f�8������4D��x�;2��-&��O�B��vL3D�z��=e&�ΐ=1��=�g�1D�x[�M� 4X�HM�y�تGK/D��ť�$����KЗ$6�4C4�-D�ȈEbXO�nx�rb�70�P}p��+D�\�B�4=t�ڄD�!/�QaL,D�83�[� M��c�,)���o$D���(� '戹4��%b��e�?D��R�@�A7�E;�Q-؀���"D����C�ZT���h�;g|�D�v�>D�̺��@�u;�Α:.��c�=D�$	�o��O��9{E��5�l�)(D�0���!(��r���7h�MpR�!D�0�M�2PY"m�*Z5M閍�b,D��葤�� �TaB� +���ړ�(D��3�Lۗ�"��P|xuB�g'D����N´s����N�S9�I�B$D��CO�3j�Ba����,H��rE!D�D�Q"�w�>a1��u���t�>D�Z�E/T�8u��(�$t.$IZuo:D�vj���)p��W6^��;��#D��B%.��T-.�Y���L\�$ņ!D��0mԕKn���e��(ĺ����?D�PR�!զ�=c��0
��*B�=D����h�pAA�+��.�t�d�7D��µ-��1���0�[7�l:6�3D��a�N��V�1z��G:f�,QAb5D�ܙ$ٶ_�}���F5@����3�2D��C�:�"��)�f��n/D�� �8 �Ik�*Qs!�#ZB؉e"Ox�Be>;gFu����*=4�D"O0HѲ�L�5�A�wd��5T� �U"O�p�iQb�~<���lG�qx�"O4 0#y[��R�;Ѧ��"Or�c'���q5~ͨ&$��m�t��"O�=��$E)a	�k�#�  ���0�"OJ��c�
K���B�;lv�8#"Op$�	��pF8�p�X[�Y��"O`�z�ט3��ٓB���8�r"Ol�q� �����˄C���&�#C"O(�6�-���BM�Dx��"O�A�ҙA�p�S&�J�2���"Ox=��ڰ$x���-��!�"O�Y�LC-Lw��A�Ss�"O�\ ��2Lu�0�-�	 �"O2,�#�):}�x��m��X8��"O�(@EY����f�?�99�"O�\�E�G/	L�#�Y�t 
� #"O����D�x�б���O�9c"O��Wo�)%��*�� �5��"O��tE�����*aiX�k�4p�"O�]��H�T)@����Y�"O�� ��X0��`�%G��T����T"O>3�,��a\���ve�W�`H�"O|9*�kԓn{���3E	*wB"���"OZ�81J�o���!e��R3L�ʐ"O��Ռ�hPũ���2�2�Iw"O�pC ��w;^�Ԍ��\���*"Ox�1�jS.�x�_�k�����"O�@�K@$^�2iI��H�T+؁�"OxT��D�JB��ƍ٤D#|D�"O����"}) �!w�@�b�,��"O�+�nL�d�h�8J�I��-�b"O�q:��ϒ9����&U�	��-�6"O��0��9����fF�Q�P���"O��``�n�B�	p�8�Y�"O�y��hFF湣��ڰ�n�c�"Oh�HIPT��e)Zq�~�!"O�}���6��H����C�"O���� tZ�0a��ͬv��""O^�3q��	����ϲm��A#"Ov���B����iQ�V�[n�=�"Onx��߳i�t�̅F]<	�f"Of���d��� H#DǇ7�*�5"OBm�W�K���M�t�Z=_�d�0"O�q3�/@A�<��`c���,�y�h�d@��V���bC@����	�yR�ͩ~��1�!US�C��>�y�k��L^L1���C|�t��A(�yb푙/{d���mǄl��pщ֨�y©&gb��X%K�T
�*@�^+�yU�K�buX�	�*N<B��ҡI�y"�L9xx�IQ���A^n�h�lF	�yRض&������3@K�L�3�S-�yBϒ��h� ��2������y2D�)�T�u�.B�F01Ħ��y2N�7�,�`#�##Sz���f���yb@_�&�s�ι �i�i<�y�	�[ATY��[�eb��:$����yR�
DL,��S
�;^�ԁ)a^9�y�C��J���qsز�|�TÐ2�yBT It8����X�(�J����y�V��T����� x�,(��!ڪ�y
� �j�e�OD�K���/��$��"O܍c��g��u�T�Y�Q��̘�"O䐠��"�ca)2����3"O�5:%�]�.�	����B��{T"O��Ys!� Z2��3/��4�,)�"O�����)-�q�.F I�v�Z�"O`u���¯h�<\�n� o�d�0"O�;�@=Aۢn��U\y7"O��h�eҠ��Ңզf^>�A�"O�h(��j���0ߣR[V��"O���-̦�	���JL�̐�"O�4�0	j�  a����D6�T"O,p����:}J\!�mM(NS�]0�"O�� ",�
5�`��]�i[� T"O`�5&�Y`�`0�0
!~� C"OT��PaF19�鋀 T�>�1��"O��C� U��4�0fS�K�Ț�"O&D)$n]�VR$<pe�HeE8Ȁ�"OҤa&��!���ʷ�4'^�i "O�(�̆��d���74Eb�Ӳ"O܍���N/(��@��l��n.�4�'"O6d��Ř�{F��E��DØISb"O�\#�0p��c�����p"Oj�)e'�p�j���q���F"O��+�A�?2	0L�v?D�di�1"O(���P�qy��8��I�|�,�#�"O� c�kB�#�����̮eB�6"OF@9L�5��Q(�$M^�M"O�p���<E��ڰፃ[[��AD"O.Hʣ��8RY�왆!OJU��x�"OP��a�RB=(� Р��� 4��"O��-��Q�d!"�ҤE*���"Oh}���*H.��'��!e�hy�"OY��"^�Zԩ��S�	nq�"OfE���
b���D�=
�HAp"O~Q@Wa� Q4@��
{�'"O�1#��Jx���&L��	��- "O�����7ي�y"���$��"OxѠG��L�����0�i�"O֘��70f�QfI͞|�x���"O��v �/k8e���#+�di�"OL��`�ӌ�ș�j�0���� "O8�KUk�+RL.v�z���"O�ᚲ�4"������s�n%�"O�L�D��A�1x2LE���b�"OҤ��g4T��T��C\h���"O��봮c
����[�SKn(�"O�1�S��%$i脩�� EEꌛ�"O>$���*8���M6l-�q+�"O(�3a%K�U��Q����4z�"O%�#l�
b"jm�e��.L�"OpH��*%�����7���y"Û���� V�L�3N �
����y�N��A�x�����$YU��z�m��yR��0M�*�N��F���F�L��y�R ����H)7�Y�O��y"���1�Z�㪛/*�vHՏ�y�ѻ�J�)�
Y3��y�@?Z�Л�Oޏo3f�S����y���'��3�揽�n �S$���y2F^�i�J���6��0���l�<9"�wH���e��H'��Kk�<1�8��}�rS��x� e�d�<Ѣ&C8g#����dT�`%�x�Q&DF�<� ��"jV�Ww*�Juşj�pԚ�"O�H1�l�
2��9��,�"(��"O�9���Q�~ ���	]Tȝ�"OB��'C3��ra�{�A�6"O$��g'Z>w2�ʸp,=��"O���r�ӢY�@ pS/�h�x1@4"O�4�FƢ�4t:q�W<�(xs"O8=����
�ջ3�I� �&h�"Oaہ�2�.��J��U���!g"O��cd�bl�);W`��7�4�"O�*L�yN��.5Gx�L;a"O�B"(ْ9���8<��;"O�$��.U
A�0�x��J#>�*�"OrTsb �  �   h   Ĵ���	��ZHJf)G�5u��(3��H��R�
O�ظ2a$?�K&��;۴%`�F#�M6&�ׂ�g�`y�C�%&B6m�禡b�4n������'����<��@b�\�ٞ��0�J�E�O�du�O���:��B�m��+@ �D���6��g!gy��H�]���݃����n#>�*����D�k0v���X��䘩 gE�Z,0����I<��ܟL;�! %�Db��sF�R*�ʓ+]�_��
p�VV3�u���m~2d#`�s����g�S���'�rq"�(:P`�dFB;#�HL�O�Q"v���(O2�YH>��%�?�6!�խ%s�d������<�'�,� �z"<1 `56|`xH��UU%����%GR�����3uh�I!�V���c�'5��=�Ci@�J��'��ADx��Bܓ�������L1���3#�Fyp�l�-������	4qH�� �/I* [�3�݈Er�xEC/�I#6���i4��P��Y�KN���^��$�Տ�<��<uX�pb�I��H��"�LN����l�vd��3�IV����69F1�0)��xll �C���'�l�Dx�`Rr�	� ��E��I9L-�8�-û	Z@��0���Z�x�^�Ԛ�N��Bep�x"M�0-&l*���O�(1t�G�<�-
6��oZV��Y?Y��, ��,Pn��U%`p�M�1.љ*�P0/O��ە I�K�'{4Ћv�ɾ��8Q��H�L��2f$a���6#����f��bɦq$��Sӌ��bԔc�ăca;���i�J߃)�D�ݯ9�v��;�fy  @�?���Y��O���d�� ��6.�t�Ջ+0 �0P�Bi4��ē��mM�T�O�|z��lz=�W�'�r�'�R�'�P�2u ie]P�ka�B�Y&�'<B�'�N��!_���	�E������
��&��'B�Y���R�5��q��� �'�'��/V��Mk�'�-�,Np�xgI��sl���ѮN�uўD��>L[�T���:f���"[-��듶y��1	,���H��v	�v��I�E�JqKr}�� �O>���O��$�O�˓�?y*���]Od�5P��1/6���?q�&�dQ��9�޴m ��	|ӌ�D���Y�޴,!�VO}ӆ���3h�ܻi:2���Q6!�:)ov�=���0r���D�z�� �W)V�wܒ �Wa/F�lAgHU0u�ҀnZ �M�i$��՟�i��ۄm̔TR��!���� ^9/�d�3׼i��]+d�9t� �g S�sn�E��ؽ@�Zc�!`�<en�!�M�w C,����HT8'�p���@jAr`	o,8��\9��6�a��l���mrT���S�d,yp�H81
�( ؍�C�S�GvF}`7%إ#���"��286:5qܴ{���hӬE9�nK�!�<p�;D��I�E�(M�T���bU, ) Љ��
�܌n��u�Tl��n>:���i!*�	Q4`	��^�� ڀ�	�1N�ёJ�.y�e�����'���'��=قuӶ�d�OXyR�"��?+��"֊Ɔ|�h�@���O����9D�p�$�O��S[�f>�aa�P����`��]�4�����E{�=O�h#ܴ.(���1�/��$���b�Y��F���6���@�axRc�
�?Q���DB=t>��r����0�� � ��'�b���Q��� �\#�<�	b���h�^���#�l�8r�� �+Գh5���q��O�D���&�'�y%F	������ ��V�Ԝ�y��2�d()�C���)��2�y� X�N��H���z����s� �y�A�LdFz�d@^ �s��y��=�j�@��7�����+
�y��(�q��*5)��+#�
�?yՀ�~���������(���J�f����$�(D��oئ18(�B��`%Y�D'D���f/i
�c`H֨b�0a� D�h��Խt��za��<q~��F$D���W*E���a5��MӚ��׌6D� �C	C��}�F��f�a�ɿ<q��g8�$g�������%%gI.9�H1D���$%��y*�H�e��3�*�X�C*D�D�RB�G�ݛÃ�0��� p	(D����G�0,���)A�d����%&D���D�6��w&�; �n�hϓھ�����V&3�4���d�!sYb�2%e� #ax����L�jM09�(���]��|f��|%�|�U!�"پd�����@YT-Ey�@	EQ�0F畺2�r��L#s+�cdlE>\��D�	���A����8g���Dy��H��?�d�i!l7��O�yRꌻ�
xH�Bэ4*�8ѫ�O����O|�d�ON��:c�PsP����>�*S��|Z�e�$1�O��	,8N��p��%'�L������d;�	¦z�(6��O��ݨ'|qa2aB�g4 7a-{B�I�k+�,�@[�.��]�'�Y#�B�I�Ul
	�g���ʐ	BD�V4�C�	/K%��ф�O�2(�2�;R��C䉶�]/�Jl�#�C�4���"O:̉#��k����.Ĵ8ՠe!��c�l��On�dͳ�th$��O���O����b�h%��K�9���l>U��a�FJ���""@ɦ���f�?_�zP�Oo��xsdΗ$�bU0u���)+ Ź��?v���sB�z���A$��+2�c>c�d��h��Ե7o��3n�܉ ��O�@�'�ʸ��bY����'��tg7o�nY�>}�x�@֯��"O: @Wf#'�~Y�bN��\���X�� �4���|�O��$\�E�!L�z��	��T�ht+2�I")�:�)��W����d�I�?���쟈�'�ҡ�aL7Y �`�G J0=����&��Ȣ�@?Ohp���kмZ����pc[H�I��[
Ɯ�N�����	�z!��q�����4�ME��L4��4L$ɔ��'oS8iB�yp0�'����~�'`�Pp��-�x�i�*x�
�'j�hV��.?�*�p�咹f��H�I>�u�i�BR�d�i�,��i�O���ANNjٜ�	��?!(���#G�O��DO�L�$�Ot�S�]��<��&1ePe� �Jҟ� ^�S��4�r�9 �"�����'p�u fm��/9P�醂;��_�4���P����Y��ӳ�0<��OD��H�If~�љhrl���@9�j8�����0>��M�U�X�`���@���p��a���a��`b`����19���	�JPN ��Ixy��/F?r�'��_>5�m������)�+>L>�r1��*m �dȟ8�	,?���s�Vk���L��
�ߟ4�'9���[�+��`G=}t:<Ir�=?Y2��M���I��ˢ	�Eb��
:��r���)�<����e�!ZdLûb'�"ѝ��[���O*��=�'�y��s��}Z��M�^Tb�P� �yb���<��8�$�Z<,�L<B�'�:��OiD�t��/WzH�!d�K��A���I6�V�'R�'n��grT��'[��'���^�|�BC��=1����_�1OTY�R�''"�#�J:|���i�%���f z�y�����0=q�����w�q7��i��[̓r3����T��Sɛ�Js�2��Pl�zsG$D����T��e{�I��+D�h�	��HO�I/��ZT�}�G��jc���"ڿ'S�A{` L  G<���O����O�y�;�?�����$IO�_�f��	�L��x�jF�f�hw�J-� -��L�� ��yRn��,��T�&�!z�s��M�~2�IÙ 
R�����0=��ጔ����Ej�Jd�կ��N>���ٟT%����۟�?1�a��8���I�l�;|N ���С�y���&R\�usU��VW$I���X��)����'A剴;�DI�O ���P�"D�Q�@�k혠�ʆS=��$�O"����Ov��`>U�"��t�\|%�� ƤULH
	9I�3jS�5�q�:O
�{!�D�H�r�O�uqۙV�DBC�ւ-���SB�'�̴���?���?WKɐG��T��^%�m �b����OZ㟢|���9+�i��H0{��M;�l�R���B�{�(�Xd�G�lC<(�g- JX���PyR#Ũ9��ꓵ?)/�@!3�
�O|�b�唘.�4qKW�ߐQ�r�"�n�O��Dѣ@��d�7[�g#U���'����8E���h�C�
վ}�a�_8S��I,!IN���&��I�5s4.]B�O� )� �BQ��Kg���
g�[~ŏ��?!��?9������ׅA�]��E`�T��\��&�|��'�azr]A�f�
P]�R�f�Z��V9��O�\Dz�ك	�hq���Ly8�2gA
�F%beɘvJ�O�剟\
�`�r�އy���۲��"H#D�@�P�
Ax(xq��K)��9p�+D� A7���!_j�j��M����-D�ē�
Du����V$`E�A�B*D�X��*[�O��Paψ�m=�*��#D��nT�o�fT��,�a��1˓�<a��M8�*��!Gb���ǒPh؁ f D�@7�[�L`p0aQJl��[E�=D�8#��O'U���p�\�8dTQ�4�1D�\I�MU�A{�Ԓ7�M6(��%yDf3D���%&還�ю�0
5+�#�O����O�5��Q�&�V��E�5ZgRA��"O�����*ID�Q#�	�\?�<�g"O���H�)i���7��r.�ЃF"O��ӣď�{�5m:���P"Oph�u,���8��Pc[�%��"O�	`!��@Y��3�a�)zr����I���~�r�D�b.^�c�ŋ
D<�y��k�<��	���{��y�!��f�<��ԌV�e�Rk�?x1Ne	 ,a�<ɀ�Ɩ)�aK�I�����p�f^b�<�Ǡ"l�`�ʠD�1Iq�L���H�<�4��;8�r٨�IQ�z� �c�KO��@x��(�S�O�d9���#��%��X��B"O�lk�J�CʒLb�oW<`���BT"O2ȣ�S�Ba��-8:T:d"O ,�!��}�����uS�"O�#�*lE�x��ڇ���!"O����ē	n��a$�J�<�2l��_�D*�i.�Oj�Ɂ��|��8q6"R2?vdJ "O� ��Y�.k~!9�̙wQ�
�"O�mr����3)TŨV@��#�"M�"O]���) Jh�H4/�}�<��"OH=�
[�dCRx��W�-p�s��'�f���'�>x��ۊN�F���N-��a	�'��9�E�b_^� �C݀Wݸ`��'C�E�ɌDv80��GU&@�L���'o��X�����$��nO�C��հ�'$��R)�Y�� ���(7�f�{�'�h�pd/��t����7�Ѹ(-�X3��$��e�Q?��E
+>���kn)<�rk��$D�|�dL�6����E�P�,8�`-D����˞%	B�3��O�3��0٠�6D�����cPDIqa��W���6D�<0�Dba֋I�7�x�����Ox�B�I�jS�8�l��L�N�j��ܕXg��d�?l6�"~��]�O^~9��1PNM0�	֞�yR��3p���Q�� �L:fA2� �y������)��VC)���'>�yRc_8|����*@��e�&���y�آYb��UL,!���2u�A�yҁ�C(���P�"��CWcŊ��$����|JC�B٪�hϦ��̂G��0��[�N2�
ݰZp�4�Z7G@��������MV�_^���2o��.8�݆ȓ$��1�֓;�t����/��m��.�`Q)c�ںfv������mvn�������ɻ���G�J�$��<Xv�VRB��9>�И���M�x�ִ� �
.]�C�	�ZM�4±IY;-7\I	����g>�C�	�>�č A�ŢW���"��,��C�ɦZq���D���{���`%�	�x C��!M�n��BkNt��])�%C:}��=����K�O�t
� f,hB�,q�����'���YR� )�<��a�n���'������	��@8q�T<^� �K�'^:�+�ʄ3�D�Q %�e�~��	�'��P�d��.S_V��J��T�~=��'��Q�G���i���GԂ=�>���Ex��iлI�� 7�9��E�R-�B�ɍ>�֜
G��y+H�JEA�SnJC䉱a�������.�7�L*iZC�Ie�`���ٚE/J�X4	 c{�B�ɇ��`�6�X7Iޭ�$J-I�B�I�P®��p��gqƵ!gH��k5<˓G`8��	�n��uⳎ�0���ӃB�Ob,C䉰-` %
D䐙h�4�Ѕ��*C�uP�p�4��%r�Z9"���w�B�	67�����j�l�*���T�LG�B�	.XfU#'C�5^ì�ʦᑤL ���N3��D��n��D�B�	p���	<o�!�d�2'��P��SBT �P#P� �!�Ѥpo��K��^�(���7�!򤒗�8�z��S+8��X����!�ή#�����@�9zz�4)1)�j�!�#e焸Ǭ�8i�h�3e$wў �4�&�'��S�ݳr��xy��k�����*��5���( ��M
4k��ɇ�Q�>���]|.�	ñ.�0U����(���`%���AAF�(A�ȓ'�:�"����s,6�X�}Js"O�$���16��X�lءs��}���'Tᘌ��ӻ
F 0 �Ö�J��R,�p��&���;�A�Gf,��
ԾV��X��S�? ƴ���?5��\���,��u�p"O$��W��Mh�JL��:�J<K�"O� �� ����P7k�,�h��"Oy#¢��g��ؓs�A�(Ղ�ےR��ɔ�1�OΤ�f��� ��Gʎ��"O���ՇʶC,p!�z̋T*O ӡ�U�	�P�G��VT(�	�'0�	s�`��5c�tIG��:��Y��'�<��!��/I
X�F`�!,tn]B�S�����a@�@�*�"a��1�V-��8۸$�B�\,�#)��"	�9�ȓ<|	s�c�4_����N���ȓT���C�� 9O0U�!I�)"��i�ȓ	�� $	�X���M�(����F����Û�Uܘ�6 ��؅G{�a�֨�������q�l�a(��&p�"Od�`��ro4� @�E�pm�ِ"Opa��9��%8B)?|UB�"O6�ӌ����ū�-�i7���#"O���g�I6BvD`L؞m}����"O�9�hfP!�vAGu�1�'p������#mOF�ȣ�I�J��(hR盜/h�����iV �:I{b�2;��B��;(���k�u��`[ 3
��B�I�9Cf\Z k�=s���e靰-fB�	��r�{��[PNȹ���I`VB��7nS务��'��8��n�'�Lʓ4`����# U��Ń�';	+Ԃ׎_�"B�	3&�`�3�߄m���j��(�@C�I�(;�;���.!Iƴ���ߏ9��C�I�Kj@��	B�[�^��n����C�
�r���O%l�y�#W�c1���Ĉ8����;M$���-,TĶ���ы�!� ��r|1�O^�kV2��v��Y�!���3^�v��ѥL*!�� c���!�DĈ"�<m�#�Ƶ8�$<z��Q�~T!�dZ���9��n�V�\,s"��qr!�
�� Ց�e����@�pK;E�ўP��:�C�V�����P(�en+�@C�	=1gH ���7k��ЪW#Hu�C�	�'�L1ॆ�_���Q$d�w��C�Ʌ1�����Ή@���rDI"R�C䉾qT��q0�@�vl�`[���3�HC�I��)1wIW�Q.��7��^��dD�h�"~�(N?KÒ`�rÐt
��R쓘�ynoԾ9�&�H�7<4 �Ż�y�e׿#"80��m�2���Ufф�y"D]O!,(���X8Nb���̐��yB�<9����I�f��d$R+�y�(ȮS�:)q�B�\�Jh;$����$�>o�|�!�NK���a�C���a��V��y�+Z� �i0iX�h�|��"!��y",�êUۂF�1d�r�9�y���d���0����a�)�(�y���Fk��a ��
��#CΣ��>1Ԭ\?��ȐV�$)��GI�X͜�I�J�<�6� �Đ���.&���JE�<	W �*vw���.�}�\d��eH�<��I�q�v�FJF�$�V��e�C�<Y1���j�5��O�V^¥��|�<	5d�f,\ #�\��x�!g\B�'����iCJ
���a��&\��I+A.2�!�dA�BT�����2xp=�����!�dD-J1�q�ͻsl*Z��=�!�� �Tk���'%%e ��y뤝�"O^4�V-�$�pQH�$�N͘4XT"O�LX�!���=��@Y/b^���'�|�����yR5����8�E��N+ I��X2&�C���}F�R�}d>`�ȓ��=A���B��� ��S!h��ȓ8Ѡ�:�[4w $��ߨ#�Ԩ�'-�qG,=:9d� ��E!"6�uS�'�~���l'?�v�Ka䅼b��+OA ��'�ʕ��$� ��q�3=��1�'9�A�#	�Ve�%��\�m�%��'��<A%ܠb����c�q`���'����I���Ɯ�D�@;z�'RT��cI�<��u!�I��p"> ������j��7"@=��)���/�̅ȓ8z�[�C^�s2ڽy��6Z`���p�g��TN�A+�d_.��g��'%�>�Rŉk�hM��
�^�H�!�7k'F�j�BG�$()��o������!�dR������E{2��˨� ��)�!��@y���;��"O�S�)>������ST��Y�"O�]�'�՚hl$U!G���,���A"O�L���i�tȂ��\�_ò�*"O, Jŧ�O�`,���Q�TLJQh�"O�h��	2H�D�8JL�H4r3�'�b�x���S�!��щ�e�5 B2��G�����>�rW�;Z{� ��2�v0��.���&��%b�v&݇E�.E�ȓ,��HqF�B�P����]JN�E�ȓD��1���HȖ}�Gڻkj���Ɠ1P�[��8����(Q1 �@hȋ{��ؐ��$F<vy��'�ҙO9�TB�#� vfbm{�M�
$.�8��^&\����?A��"i0����I "Y�2k�>ͧY��T �HȅU�y������D|2N]>Oĉ��X�>���t����T��š�C� [\Q�2��/R����Ob>�� $�p֎���.��gD�<	���=)Ć@l����.��5�����I��)Ĳx����{�����R��9��Iޟh��O��R%e�
	簥b��Ф2GDy�3O61���16���Ba��o}��I�#�.�۳�]�J��C�L��"<������.M�2�,է��Nu%��<	f�P�gʁ(���0�;O ����'Or����f�~�	X�j�xe��Y!��$T�ȓ���Pc�nݪ��鉴!��eF{b�9�'u�"l�����N�j�'�]��Բ���?a��E�^J"O�-�?����?������)48{PO��c�|swL@�������Ω0�TՉ���V&.����̟f��>IAr���҈D�#&��d��'�ٗD�(�6`�$õ+O�8`�?ѱ�4�M�R�������L�:�)Sc1)���K��*?ic��֟���Y�'d�½h���s�T�qF2��¢��mD!���!X���פX0Ѻ�ȑa�=�"��|b����D���r	�@��&%�#H�"6��y� �OC(�	ҟP�	؟���Ɵ`�	�|��W�v�RԙvmQ��Q�Ūs޺	��Z�&V܇f���B�	s��h�4K� q&́z�)�n\Tr����D�fP�A���6ǅ>�Mش��O�H�'������3S����X�f�"��'�ў�F|r�J�}�t�$ ��v��k���y�΄�t�z��AoI"E>i�fD�'���¦-��pyb�5��'�?�O@`�X��8X�|�٤�ٔZ�:����ob�����?���t�D���0i�<���e��]��Ou�5�'�ٰ�fM�$ y��ȉ�Ą�?��g$Ф-��4�é�|�� ^MJiq[��:��I)w�h">�4�����	Q̧��y��Z*Bm����9����'z��'A��h��#X���z"�թHlJ���7��C����^ s�V��g�M*���q��YK��io��'���78J��	ퟠ
���=��9�q-H�)q�	�'�㟘CïԹ-�������gb�3�S���\#T�t��c��9:����F.��$�,6W���rfO ~ٴ �"0��W���F�����Ǒ��� ͓]�`������'��� ��P���-��d� ��pW����"O� 8�%�9���"��Z(@3Q�"�ȟ�(���#@v��#M���vQK��O���O��A&�I�=����Oj�$�OrU���?���6v�	�"�W?d&v��aN]�D�d�'Q�=:��J�*��� ˟�h���4�8Z�柸9����>h`��I7t 9��\9�@�g�'�h��C��[Br��`��u=B��O��*��'�b�'��O&�S �u���L/ (ЛU�t�,B�Xdh��aŵTfNqc� A� �2�d	S�����'��	�2$���AcH �ࠌ>3C��F�
_4��I�����x�SٟD�I�|B���-f�P-x�B��%p��'Je��(�'	�t���ՙxڷ�I�=*)�	ȯ	�$L�YE��Ǭ�0sִ��<I2F�P䉞3�M;ݴ��O@�kp�'E�IH"�_�V�����m*`½�G�'ў@D|R ��X8� �&`s�됡���yB�`�Q/b&�"���S��'2\7m�O ʓy~��ܘOI� dK�p�,�a��}����DC8*sh�QV�Ԛ6���S�K�!X��0�(����En���F�p�o�BG>9S�򄙩�r"I�+��q�k�{ ��R�KZ*+�J\�C.N�l���,�AGz���1��'���'D�鏻i�8;Ug�2���Bbi�l=��'A��'��R>�ExR)�af��q& .��S��+��>Y�]�x��k�GwnD���2-7�K�
�<���ߛ6�'�1��X�`��hQ ݹ�dT�ɾ�	T��~�	T�'��,p�	̵3/2Mz0L�5nr����iU�'�&5�|��	��j�������<Zv ��CHG~b����7}*��$C�N�T쫃�F�9i(�9c��;EL�q�!?�s�>!���Y�$�x�Ӵ&���"!�(פu0��
2|�]cR�>�p�O�}�4�B�2 �/1��<Zf���i?�ʕ	Do�dTq��K� A�t�S�e�@����7Sș�a��'�������wCEE�"Y��Vi��y��-`��1$e�oԆ��I9��I)V9�'�z7풳�~	�悗P�d����X�I�_��'�,#��hG���qb�Ù;�&1��ϑ;b�dM��S��'d����O �R'E�g7��ZA�=���;�c��uR`� �@��'�j���'C1��i���!�r��$�F�|����q�'����8����9O�y���O q@1�P�W
��3&AϠx�(�*��'Vi���/z�Ny �G�i=6XwCH^��C�ɝ��=
%�ްOt,h��j��&��7��O2�O�1�����|n�Q�leY6�5,�x�g�JT:��䓺hO��r��r�)��=q�턅t�.C䉀��h	Q��<v��i;0oğpC�	-uɘk3(�)+9���u!AK��B�ɿp�*E��-,_dȋcg���B�/G2F!A������@O�d�&B�	-l�,#��ޱH��i���ʬK,C���)��%�Ir��D�ȯXK C�I�=���«ٮB3|U����=�:C�	:�$�����U�X)Q��<�HC�Bxe�$t������ؒ�2C�	�_l�I�g��-�p��\>�C�I��S��ۿ�c�-�_�C��=`ޮ�+Q��z�6�)6������2��аxǬy��" k�:)c�()�4}k�M�2f�)���n�`�)*X(|)�Ý8x��ƈĘ(�Z5���?JE�,h@��Z��<�-W6@ȉC���Ik�a�!�Of� �h�&]jT�u��+z�0�	��u!�)f4R����7(�lQJ>���$i2���B��bO�R�FC��>��p�BoD�(�B�;&��?~ C�	3ˆ�@�yj"5��"�\C�B�I�?wش�+˯i�	��G��$��B�I1e�,Yp��R�4��C��,2ZB��6^�
x+a Y8@�`'��<�,B�	*.��x��鎑PH.��g�B�
XC�I�!ZJ�hsIA�&��KxC�	�B�ڠ��<��e8kH��jC�v��9sҍN̊u�s��	j\~C�ɦMC����+�8��E�[�HC䉿e�4��q$B/4zIt�D�@C䉻JD�+�*ϪQc�xt�ߎl?0C�)� |�j7�\.�qU#�'� %� "OB� AB9�y����jM��"OpAe�/	�y(ACN*N=��R"O\��w��]NЉGA�Y P�z�"O�D�4%O�A�ZP���N	<�PW"O�iJ�G@�FnT԰���3V<�P"O�,�b��h�T=���?"�����"O��b��8�.�bc߳8W`�g"O��ǭ(ղe0��ۈ ����6"OLA�7d�&m~�QBM�V�R=G"O&8��,R���I.
�5��"O����L�%�|x�6'��f��<�5"O�T��ހ|�����Ky�ĉ�"Ol���ȓY�L����S�.�4�"OvA�T�g�PcIݸa� B�"O~�I� �0Lz�ȵ╭KЌDu"O�hwe�b���2�x��f"OR�&Ѩ-2V� �ȥ1�ti�a"OT��V�06���!��.L���"O��{��ѠDri``��:�d\	�"OB���%:$�\y`֏��f����"O�l��M§�B@�T ��#��L'"OT���5%V�rPn��Y}6�X�"O��bzI*��(u����e"O
mArF�+<��Bb�#oh��"O>�q��Xy�����I	uh(r"O��@�����JH�^x�!u"O� s��5"���C,P)��#�"Oֹr�ʗ�Q����� �B�&<+"O4�1��sL�31` �Z:v1�r"O00;5(ޕ���@�/;4�0�0"O�|!�又}�<`��$��.�t���"O��p'յQtɠv�GK��li�"O��el��m��MЃ��+�|��3"O2���A�|v&X�B��My�iW"O��a��=�Z������<вp"On���@1����ք�V���"Ov�;�˕2ςM�1��`�(�A�"O´qB$)%��A���Y�	 �`@D"O�9)u�_������@8ؔ��"Ov��"K	�8q�U��u/��C�"O�ш�,��E��Al�v�$�"O(����A�_}L��k1�4��"Oũt� !ɪ���_%���8�"OD0��5A�P�㊏<}���"O��2��$�6�H� vF ��"O@��T���趭�5t,�i$"O���e��UK�Z�iW�u��"O�8sL�	:1��?>,u�"O��Pt��-X<UR񲢺���@�L�<1R��jH���P��,�j$��&�s�<���QIr�HO�@Ǟh�Q�Z�<q%!�8F@\����nnRd�GL^o�<� HC����D$ϻ�"��B�<�QB�V1�lӒj�1C���:��S�<�E��]ꐜ2t�G�s2�P�<�2��m��e��@�5y��r�DE�<�oD�# �}�R� ({ ����<�E�V���	'�\#�Lw�<	�)Ε]�8�@�C��L_�#��t�<١��f���"!�!u�U��X�<��ʑ��u���s�z�TM�<�E <�L���̏R����I�<1��[8�B�2�/R�PI H^�<� �a�G_�hB�E�5�X�sT�|Y�"O��C�jL�G����&-G4Z�"O|�p�O\��,���>/T��"ON4��J�>j��HC$�)`�!�"O�a)AG>D�zw�L�u�"I�"O\y����E�2i�i�0�=�"O\�9�P<��v�L�=�@�"Oֵ�e��1	I|��B`��C�m �"O�hJe��*�!��͋�e%�B�"O��C�*B�[��1��~��:`"O��B�6��Ċc�ܰ\�,� "O��K]x9�J$�$|�4�"T"O���$�6�|pH��+����6"O�I���'��)�b���up,��"O�葶
��i�Z� �̞�6c��"O��HǍGC�b�У(��Je"O�ts3$�G��rʒy���"O�0�#��(nԩT�1'��(S$"O�9�:sQ� '��$ ,m�"O�ỷ��h8ii���Yڣ"O`�D��$c�(];��KB��"O|��@�d�֩[������u"OD�ذ��j��k-v舰X2"O,�곫A��M�P ˊԘ%	�"O\�jC��_:��s��Ǧ�r|�`"OD���-�E���.�_�5Y"O�M�T����,9��@�b�5�P"O��H��!,6��Cl��c�� �"O���"'�9k*�X���ؐ��EQ"O���HM��0����Y���P�"O���b�����7@��y�C"O�4��l��8P1/�'ⅉ�"OB��TDۊF�8��`����H�"O��s��ja�Q
Y �>H�!"O�����zמeI�nZ�?���SV"O�\����!HX�pCm�F���"O�).Ӟy4�k�.Rؑ�"OJ1�aZ�nx��쁮,��(;�"O�r6�� gJp�;�LB�r�sC"O>����ڰ=�2i@"���~�S"O6$����2���`��C�9��h��"O��C�
L:a�&�R�Eڕ`�����"O�X��F�)IMN0Z4F��"��D� "O	BoR�cA<�E�V{��q"O��A��Vs���ذfD4���"O`�	�??����"C�*h�!"O&�1�<m�<���BA�t�:�pU"O�J^-@��v^-G攀т"Oa�d�D�
��$'� x��"O8�A�lUf�h9d 8xЌ��"O�Q��O�C��P�sݤpQ�"OR�H���h$�5��cڙG�}��"O�+�녤c�n�pç�+z�*qaT"Op�A�CѺQ�"aK���F�j�3"O����$t�^�0�e�,u��=*�"OFL�F��3cs�!�g/��8h~�H�"O����%̮L !qN tp��E"O�S����@���`�\�S��ī"O���ú�a�qnO��=��"O,X��1Z����&�sܬӆ"O9 0JP:$�Ԩ����$gR���"O<A�q�Pv$ �U�F��[#"O��)1ϗ�4���(DA�B�Q`"Ot�(���z�e��ز^(��"O� ��`�q�<�s�R1%�2X9�"Oii��4=rE�0M� 9jN	��"O�ز"D��e��hu�Hqc���"O�<ȁ�T�]��FkW�\EJY#�"O�A �B�'�D��S>-1�H�'"O�Y�C�x������*�;�"O�遊��8YX�`�F�n
QBF"Oܘ�5��F�
a��$�FYpt�e"O�=��㊸+���3��{O!c"Or(AL	�A+D k��R�2��8�"O�I� 	Nt�h�š�b4(�"O�,��dΆG_�EZ#-��P���Z�"O$\�$(ۨph����"�!(��c�"O�4���J��Q����a�~Q��"O�1�(�!S��B�o��xl��ʂ"O�z��Ԅ��G��-&���"O�,��#u�Z C��';�q�S"OB���!�ՙӄL�6!^��"O���vmI�3�	�uJ�be"O�C�$���l��G��3�\�Y�"O�t�%/��r�@S�d�>z�D��"O:�#@�Ѝ�&���2e^�"O2�`F@�+\xe�&�ԕ%D��"O
|�`�a(�]��Ę7Y���"OZ0a� �;jX�\J���](@���"O��sr� *�I�$萗\#|i�"O���Kʹ%J���ˤHj|�@p"O�iٶ��|J �����N�̊�"O�=��6_�@�*���U���h"OҘ���H�Ig�(�!�*n��8 "Ot�HT,��G�R�`�T���36"OHE
CkB��HB��*"��"OLQCʃ$6팀�"�L�!�aK3"O Ց�N�E5Ԣ&L̂*�F�@�"O�çI�jI��1�TV���(s"O�4�%���g0����
/�>��"O�%Ǒ���|��N%��� �"O�XP%BI�b�^)��ŀ�i�,��r"O�ĸ�-��E�"��vjگ%6��"OH���ͯ�: 
�� ɜ0�H5D�tp��Ud�x'�]�zJ`H�4D����!:�R]9� m0�`�?D���/�Q�����ߌ�X�d�)D��*1�ݣN�D0rG�!M<Y�G)D�@h�)��C=L�z��;eh����(D�h�d�1h�]�0MX2"���A2D�l`��
5l>,B0�H����p 0D� �u
�d�RC�gF�z�����-D�,K�I�&��8�3�
I�`��*D�`�	��<���6���~&��A�;D��
¤�66�P������腐0�>D���"K��5'�E�A˝_�!��>D�4�$�ψf�DC���v��QRV�9D��#%��5���� �>e��P��:D�<X��\g��8[��B(��""=D�H{��K���b�_�K,�4y��9D�p�%GŕPp�hФ��2��H�@�:�I�^�T!V��>j.��QB�6%ր�O�͹�$U�3���T.=~���"O�d+�A�}�0$�D�#Ef4!�"O|Q{qm	7F�Ĩ�S�ʪ
E ]��"O�E��9���H���"O(1�2ˇl���r㓹va�� "O�}��"�s�����_3�Ѐw"O����� vS�m�p�H�@(3�"O� �D���C�6���A�6�-��"O>��2�F�#�[Saj�9J �X1""O<ځ
P����؁�³<߼U��"O��#׎�&Pg ��Ҁ���@"O����صRZ�a�T�L&vܠ�� "OFu�ҎÚ{#:%���Qlڄ��"O*��2c�)\�p+F�	�2t���"O0j5�':�؄Dh�e�V8�y",ٞWVrX��%A�H�๴n���y�Ș�aF3AO�y �4 ��J!�yR�C�T[@ej�.�oz�:��E��yr�W�U.(�� �;j9�pq���y�$�9A6&���C�T;������y��9��XK6g�/F�f�v�;�yd��\&U�O�4��i�o
�yR�K7],�ЁE�A�ym4�s#i���yr䚟&L25Xp��5uF�� �¬�y"�V��^�r�GDE�����&���y�O9�$m9楁=vO�A�D%֢�ybK��Qz%�V�v��1��I��y��φ+B�m�'��m�v�2����yB���_�f=�AjQ�h����nɧ�y�$� vP��1.ń8t�l2 ����y�`���ZhԀQ���aڀ���y"I�)j\b����a0W��`�C��"n,�A
gH*P�j8 1Ι�0�B�	:9( � �^77:@�r�.�B�IN�1Ѷ�.t%,��5S�d�B�	!H�� :���;T�X=�%��57��B�	QV(|�B�
nKrܑ0�[�<�B�I�:VV�� Ub���';8���m�j���`�.^�3`�`	�'����`F�a���c�_��d��'�,Ȱ��~"��׏�=�M1�'^8u{5m�#�9����L�l5q�'Vd�QłD�0��5DE*7(��
�'aTM��!A^~R�U�9�*��'���kq�N)�F�z���&%��"O�d�Cm��mV�����
c&f$HV"O����!}~0�çGK�c|0Hq"O$�e��2���9����N��Z�"O�y�W�A�����
�!�~��c"O4q��Lqo��#�i�jg�}��"O~�ط��;����T���S�ΜJ�"O>H�e��',I����V����"O͉���gh܅���$�gf8B�I�'sL0�!*�tQ���U��PC�IA���  ��J����O���B��.vu� h1U� ��.N�=�C䉹/��� ӯ_,4��%)!���C�#,��(�.��1Ȥh4�L3�C�	6;��I� ͯR����Q��.wjC��){��@��9-b)3̐7!*C��

E�X��b�5�����o݁uԴC�I�Pub�.HwM|�����C�I�
�\��� �x[<@h4�ҿE0�C��&w&|�Ă�4;4�"�(�RC䉉L	FH���U����R�^��C�I�%�v@s�	U�=Μ���:l�dB�I4��)b`���N����ɪ`��C�I�PB�A�kH��:A�A㖯P=FB�-#@�
u�IM$����;p<B�	�VNdP�t�	$t�.]* n�=B��|���h��P�TPJ��	�� B�)� ��9r�64ȸa{f��%Hċ�"O�M��-Ԋ:��lyp!ۺU�b�K "O�b�E�m��9���2ϖ���"O���ȺsZt���ͽ,de��"O>��AIM%��#SN�y��x�D"O�`�u�U¤�2�BB/wN����"O$�b@�<%'`5�w˿%����"OЌ�N�4 �.�R�M�/?,���"Ol &�L�Cz�jvm�Dc���"OJ�+���z�f ��4P�1��"O���P�s����3b�2��с"O$
�a��P���@���P��q"O(T�E���)�� �*U��Q�"O�9i�<��(����!�beB�"O�	6�/xm�c��+:��8"O����Q�nn��0%I>�JAps"O�lڣIׇFI�e8@�Z.��u��"O��سŔL�X��PlI:f90�"O��2�׊
>0��',F�H*I��"O�օG-����� Ė3�:�Z""O���*ɧ9Kڐb3Ac2��"�"O>kVfT�_謄�"��Q$��{�"O*� %N�D�p��zx`�"O��0��.!M�%��=)�R;�"O�����ҀK�L))�"ќqa"O�8��hɅN�|p(q L�H�AP"O(r!�Z=Q˜dxէ�=^�Y��"O����	���5`]�6��g"Op��ʢ.��hA����
y�Q�"O
Ik`ϥ\K���V�wR��"O����S11�D  ɍ�4z�Q�2"O~����d�V�Q�����j"OҤ��L �h�ɣ�ꑸ4�FMh�'~Yq7�6������WZ��Y�'O84� ��$$z��[�_<T���2
�'!^�j2�����аu�҉��'�RQ@T-ܣ�W=oF�`�'U�(uc@�za��DȚk�r�H�'N�;cKiNfa����e;p��'��尐AAj$����H��c�'����Âܑ]�T0��U/^��A�'�h�M�,~���X��73��X
�'cι�ZhĢ�J+y�h�ȳ���yB
m����&��m�S���y�N;4��Z�h(&��(3��.�y����H���!�&]��g���y��P8��e�G��Jt΋;)�,C�ɺpk�p�A�!#�`���-�:GBC剳=�\s2�ȨI����+|�!�䝜ph�#��àX�P� �j�@�!��B����46�=*��Nx�!򄂦S/�����<!:5qC�z�+�'Pcw
��R�6�Sb�8L4���
�'�Zͳ�C�s��r��&`��	�'q~�	��^2g2�Y�+:�Ќ!
�'�x 7ުz�<��0 E�<�@�K�'�``i��[�#CMB�CĐ53�%��'�����KL{ �{T�V�4�"!��'Q���*	�]���*��2
�'4�icsFC0z�>%���84� ���'�T(`��<*$���A2V����	�'Ϫ��ā\+y�Fh�`��Thت�'�PZ��D;T�A� m����
�'��0s�˓�2�a�'I�![?>��
��� ���Av0���j�%�"OB貤��XߠQ�a�ށ�r-�""O.8��"NA�y(��w�tJ"O��! O>��u"V�DU�5P�"O��Y�8� ���p���"O�a3脬�0��7M�"D
�"Ov5��W�j�lQ�rA�^��q��"O�\9�i�8j@�:ǭ�Q�0��u"O�IH��53��0⣂���d�w"O졲�IǓ��s"L�9�hh�"OR5��Ě%hʄ��A!`��|*%"OZHL��l�r�����"OeU ��.@Lx;S�ג5>����"O�����u"����N����;�"O�IKS���i���j�
��u"O�,����r���1�d�455z�3"O��sB���X��8��E�s>�b�"O�UӒi��nE��"!`�>
��{�"O�0 ��*	[��s�'�4��!w"O搑�hD�{�z��Qmضz����"O,<�F��714��ЬP���H�"O�ٰϔ�\`䝳�c
�O�^iK"O�×��,mh⍳��Z>���A"O�c �L&}�Tc�Ŗ
�2D+"O�DKSC��T�`k!G�։��"O�	#/�:$z�̨��%be�i"'"O2@P�è<A���ui��"Od�lR�N<�ēF�ݎo@����"O�����H�������@"O�=���ר_3�
��
{�����"Ob�j��

N@䩐=a!�{	�'�#ʙ=iK�IS��ĥP��
�'��횠�

Z�Ep0X�N~Ix�'��$Pf^'9(���| (���'��Ô�"xtl�'W-m�Z}�	�'��1�`��C���a�1]b�	�'L0�(���*�4g�;/йH�'O�����\)ab�F��v<��'��,��H&,I���L�5�L��'�� ����
������+���`	�'x�Y%%աJ�������{�f� �'�P�zjÈ)�i�Wo؄t���h�'��<�HM��r����f�B�k�'���	���8HDh(�p�A.`���	�'P��ĉG�"Nh������'Dn|y�)�:���VJ�{ �'o\(1����2��U@Ճdz�K�'=���@ ����������V���']JM��@�r��9�*�	9���
�'� ;��G3B깪0J՜y�D��'^z�������~AA�G 82`R�'���Q��-@���s���>+��(�'AD�5��b@��g*)t���B�'�E`�霼M�u�&I.�`A:�'��ds�k��i5����B���$tR
�'�TyР�D�j�ȧϚ�!LY�'r\��#��D����G�?�\1	�'p���V�J���@�2P��	�'�P���?|�>�� G1Ib5��'K�y����&hI� x��>.�0�'<VM��eF�fY��* G�^BŚ�{�����M�n�=sB5ʰ�_��a���z%�LENݨ1'��}b��ȓ��}�t�� ���Ŕt��p�ȓt�(1ا�ǖ1�� �.aL���S�? �@���+(�1��.eD�L�v"O��¥�n�Hm q-D�u+�X�"O��*ޓV�I���%_,��e"O,����*Irl)"c�I���b"O�}�siy.��GAy�\)�D"O�IJ�� o��Ɂ`���Y�\M��"O��#�ׄnX�#fG×�D��"O`i�fS#)��kƃIl�u"O �I��	�j�*��A�Iz���"O�;EI?R�U0�)�+�u��"OXD��Ivo���A)�y���U"OFQ���Th)"x-iz
��� Q��y��5.��Q�_�I:��c ��yR��6 �Z�R��I�n���S����yB�%�0���(�T��2E��y��a���@�&R	i���Y�yBDQ�q� �K��5Qcv ��y��ޤW*����i-W 9�c�8�y"�H��X�"&��LHDHZ2l���yI>\�d!囔U�P��.C��ybc֎��djg"�O�n���ԛ�y�ㇵV񎰃����Kj,e�vK�y�`A2Lw��YP���#�9s&��8�y�KK�EzZ������eb�8�y�͗��]8���	��'j̆�y"��y���a4�}>1H6# ��y�拞�حc�G�% S��;1�ۜ�y2d�:`%8���֊e��⟴�y �	�ejSB�E��{Q����y�������Wn����!1�i���y���E���7�X�j�Z��\��yrs>l�(Wg�--��ĵ�y�-���(�k�n׾����4�y��ȥb<�=���6aM�lh���yR ���b�14��Z�`�g+�B�,=�8��B�=�����,9\Z�C�	�l�]Zg���_l\�1��1W��C䉪K�&%Ô�:*���A�� b��B�	 p�t�cb=�*�����GؒB�
6���:�%��J�eK0F�PC��4GC�d E�-7�����[>C�I�!�
��H�*C��(��(HiC�ɛ( �Y!tK�~ъ���ӷC��B�I1 ����SN��B��S��0�C��1{�Ct�Q�?�2�0��9��C�ɽ�R��-@�KW$����>��C�f0��&O�3p9��Q�K��~C�2C���W�����FL��B䉖�u�V#�c+��5B�}��B�I2l$��2`��eמ1zЫĨJ�B�	9x�h	�lQ�sS�=��mD50"�B�0p�|����HO�y�uk�n��C䉢hb�+'$���ʉU�ϴ.TB�:����K�>��[e@�x�B�	<8(�����
�@ˈ��V$�J�C���&p���h6: �f,�6��C��1(���[ O*\L���lG$m�B�I�Mi1zu/Z�k��)��a��BC�<�2�j$�^�4�X5a�e��B�I�hX(���M)W��JGD�:�B�	�Y���C��2G��L�6(��V$�C�I�!~4�C7~�ð$7I��B�I%�]���K�-��4� �דY��B��n���$��R�6�I��ɜ��B�)� R� �M*%���"�gY	C3֬bf"O�t�����C�T�r&S�:,�YP�"OX- E��?v|���fοbN���"O
̸֭Ο��r�K��b�~�!�"O��cF�N
?��P��� �)s"OJ�p�k
J�ĺ�a }�4�B7"ON���i�6.��:j�'J{f�b"O���Ŕ�&�H�l��@��X6;D��� dƂ;��Ţ��6�%���7D���������a0�ΐMj�x��`3D��rł�r���͌E�P%+0D����+|E��A�B��al,D�hj� [�n�-ʆ��� �>U��5D��
�F�Bʜ�#�-6aA.D���щڣ(if��C΢Pi��T�/D�X�ӕLLj��a���3"�ِo-D�tiGl	�1f(�(S�t2��7D��A�L�u$�l�W��a�b�qm(D��2T��d�4U�WjA�}.�0��*D�@�,�~X6"�d�;;\H���3D���fk]Q�	��n_�x> p�/3D�$�sn��vL%�Q�I�s�r)T�/D�H�*�C��8ڷ���p����?D�Hsѩ��Dq�� �`��Z�"D���ԢC����B��1P4��?D���`��C�4M1�jK7y��9Pg�;D�\k�.��t���!�V]�~��g�7D�@�7m݉���6B� F0J�b6D� ˶&JEa�pQ&��_�.����4D����
0�|���ឞ}{���o?D���&�N'ʈ���l�@���>D�SS����#ٕb�B�H�>D���q�0(W�P�-Z�U��/(D��
&jџ+�u�)�.;���6`'D�K�������#��(�bL D����+K^T��M�&*��A�g"D� ��?=�*\1'D�z%���m5D�4��>->^�p�E�4Sq�c*4D����2Vlf�)2����W�2D��BE��NW���@쁓I���C�-D�\��&γ$�V�ږ�y#���+D��`��<s�������n��m3�Of�Y�$qJ�˄���$d�b�������M	F}��/A]Z=Psc/D��*�W5	B�hg��Z �b9D������Fڔ���A�,?M�]��6D�����_4c���kF�)�vŹA�2D��x���"b� Kp���,�he#�!2D��a���K��y���í�xY;P�/D���vC��&g��s�!�5G~V�k�;D���T��6���� �s�*U���<D���@��� �`a�!��J�q�S�:D��3JG�d'<�ME}� �
�h8D�����Y��=��HQ�`2���6�7D�T��[�
zɒ�7s��Y�$5D�h[�aǿD�@J�O²(�<���6D�{R���p{nT	�& ����@6D��q���ʆ���]�� mr�"1D�D�c^�$ajٹ�Z /~:[!:D��ZBl�	���A��2�V�P�5D�b�j�5���� �ɐZ0&l16�3D�ܚ�)vD�Q1��<Od���G,D�l�C˖0i��X�{�Rt�S�7D����)Rܼ4bR��K^�+G�8D��  A�$�#�l�Z�f ,��x
"O ��ِIRp�hM�M1�(��'3�����=M�Դ��c@��9�'���K����]��<p) E�'t��Х~��R#��>8��a�'��Mڷ&�N��ؑ��uBx��'�<{�%A�iu�Q��P�l����'��s�%��8��]����k^T�
�'�.U� �p̙�Dd�=c:i
�'����S�\f�$@b���'7�m�u��:Ut�)��G�g�Е�'^������=R��X*�$���'W*�[�ǃ%C+�����5��K�'M�`Ѓ9'2��y�n�&�R�'�����PZ�E&F"j`�!!
�'22�"�m��P���$_�|�	�'Z�$�P�P�p�$�KD�D3Gк-��'����Ҏ �-�|d"93J�)�'@N���@O%F8H#��+%@de�'�Y��Y�<�й��kL U��B.Y��C�#K{����bG�T�ȓ6;ڜ'�`�ȤO�#@��І�U��jg,�A�d�%a�w�8��ȓ&���5�ѻ�|�t�ϹAژ��ȓ�:)�f㖁'F< q2��ko����S)�U��d��u5fxJC�X X�4C�	3T)���"'˂R�`���	�2��B�	�	�m(�ȑZ0|Y�G�i�4B�	�X�RE���AP(�|W2B�	u*�
�U5�l����=B�Ɍ"ɰ�A�*_�q0���T��C�	�N���1���7��1���)��B�=C1�i���.�H��rdԶ�B䉖p�=`��gG�T{#�֔xJ�C䉈v0�$`�$Yc�D�a,��2�B䉿JӠ�І
KrL�4A��v�zB�I�`/�b�E�*:fV��?��{�"O��P�ަ����GBP01�F���"OR����(X6L����vo��X7"O�=�WM����S���qg-�"O~��BP;'.�M�F�%yOJ�g"OB��t����=���*=(�f"O��T�I��h��5
�ġ��"O4Q�V�]�z~����ڭn��z5"O��̶��(g͜�W���� "O�!���%l
�5(�Aȏh� !!g"O~XzB��' ���C�'��� "OY�,�J��ЂV�ŜR�<e��"Oԩ
���}/&�qB`�/Zy�W"OFdj3	�g%  .L/S$�dɀ"OP�2�D�yiHzӯʫ'��c�"Ot�'(
)h��2ϐ9
� ��"O��:��³u�z6�ڐz���"O��!�A�4�T�
��y���3"O�0a��� 9��I:��Ǫ[� q"O��׌��V7�3AjǸ�����"On�f�[8?�⁫�D3PY>�`"O��I#�AiR��*�&~hf��"Ov�)�-��Xd#dS6SM
]("OT5	0�X�v(�D��.K7^��"O,9B�"��L�H�m�\3|	��"O�p���W�kax ��ο?3���e"O��K�e��1B�����;+�ta"O���2�	9F�
�;�h��\��0y""O� B�R�
܁l�P�ٶƇ�H�ށhg"Oh��W$9�}
�Bo�BT�"O�P�@(4�>\����%{4�5X�"O��`CD_:e���tGԞR,�ju"O�@�'�=թPGI�$qk�"O����-]�R�8�F a�I �"O6y1f�I
A+2���N�J@'"O�!�%Cm00cE>G�4��"O�%ZB�¬mqz,: �Sm2�'"OL��e�Z
C� 9���J��v�s�"Ol�����^��0�hZ�}�.�z�"O�U
����4PҨ�	]��� t"O��4G�U�\ s.���tsE"Or��d��2��MU�n�����"O����DҶ,'�Y�'��QE����"O��#"�PnZ���Bڇ,�,X�"O2 �2�ܚ�:H�����4~!Z�"Oh�ʔD�
�Fp�T�8��"O�vϝ� @��U�0u,��t"ORV�U�` g&�����"O�ŐCI��4ґ�
8q����"O��@MɁ���(�bɴb�j���"OV��֠�zWl��C��!,:�$�""O�$��m�kH��g��	+(���"OҨk1i��j��d$�Q&tY8T"OL�qv�D�W�:���!2 �"O&��ŤF*Y�l�2������"O��Q�q-��3�mB��d�"OZ�r�� �
Dn�5x>^1�"O��2�L�F���r��10H�)W"O��4���T�N��E�߈/9<�R�"O�)i4aA�+���@���-��;�"O� �F.�:E6�̘�b��  ��a"O�`�����P�8u`OA�T*�)�"O�iD�Q�w8�ʡ�C�L�b��"Of�W�^:6"z�3@�6P���k�"O���� �2�X`��.���"O��!r�N�l)h$�?m#�qY4"O^���ɀ:n�`��''�,#�p��"O`	�"��9ڄYA�аVV���R"O�,QC޶X�`YSu�ã]Z�ū�"O�ݒ㢀�<>:�����yK���"O��ч^����s�ػPFl��u"O`q�$�L"����/40HR�"O������>ى���&,��"O���dіd��u��K���2"O�"�B� TP���s��y��X�"O }���']>�bE��g���[�"O&|����p��}�s#H�dy��9"O�Q��I�azh�W�I�yxn�H�"O�-HҠ.2�IЗ�P�1U�eї"O�ٸUg�38D<daPA\���"O ���3L�(��X!|���;u"O��ӗa(�����3pT���1"O��rE���z����A�ieԌy&"O�����ϫz�8�#�O[ Z��R"O
�;W�$�5+5/O�"I��"O8k���4(7�ذiZR�0�"O��"�͓!SSB��E+�<%:��"O> ��A�B�ld*E���͚c"O.Ɋ�����I�G�@5(:��"O�#��*�
 �P&؞t#^���"O\x�t���{��V	5~*���"OR��ß)6�8�qs�ZMd�Ч"O� ̥R)T�Ĩ��H� Z�BQ"O�H�&��`$�b2���Rf�02"O�=�B�`�����`D�,Lx��"O��k� ��ȱ�O�h����u"O��pa`O0/�>�+EoV�iۀ �"Of�d�j�en�x��,�"O�SS�΃[j�Z$@�!4�V�b�"O���B�)Xp�wN3 � e"O����h�=�ڵ`3-�;� �ir"OLԸ �"�|=g���=��U"�"O�y�c	���r�OX-<yj��t"O�Z"$EI�X1q�C�,V���"OkV~M��L�1Umj��u"O��q7E��s[j@�0D�/^b��"Oz�r5L�aZ�ax��^2�6Q�t"O:ĠLO�����#�(�K�"O�P֍��[��|�@�P1���J�"Oڱ�1K��b�
�N@�VT��C5"O�rDX�rX�����^6XB�"O��K�m�_�
�P�mM)7�츂"O�I��.���$ ЌW�~, �� "On�Id��u�\��K�:F,L��""ON�c��O�9ZH��)Y:C~"ܪ�"Oз�J�OĪ��y,"O��6��.t|�yQiE�?�t="O�5�4-�~��əg�Qm~X��"O�!{�h�C��Um��LTn�q3"O�u�r�� �VX5Nۦn7�8"O���ޢإSE$d ����"O6@yƩA�?�����P�%�:�r�"O��#�m�X��,1%A^�Na�"O�л���N�n	�c�0a`���"Oj�"��&}Nʨ9����c�64g"O��ug�\�9��Ƞ<�L�"O�a� ϟC�.���٩K�д��"O��PǗ)V���膱9id0"�"O�8Ȥd�(�`"��
�B{��b#"O���a�	!Y��s&FGPn�ق"O5Ʌ�Q<?m�9r�OH��0�"Op�Yt�=`�,�D�s��X�Q"Op�1/�<��c���2�a�"O�h{��
V�HT�`�41�1�"OE�]/6�G���S�"OV; n��k7h9�u/��4СX�"OFI�%O��HӺ 0�B�a�X�"O�W�A�ƭg�֐��"O�$�G�ī7�L��0�
���X�"O�f	�OL��ʒHF�JPN�
�"OP���Q�+�Z���gO�.*�83�"O ���_6,��ǲt��e"OĠ� �O*K�fX1^d4�S"O @�7mЯ�Dl�eĞ>����7"O a�Uf �dq>�O3�� �@"OQB+��s�b�{a�P���W!��= ��YibL�O�����K��VQ!�D�K���rf*R%Q<�KU��<l�!�Tj�MJ� ����JT�ŧ�!��^F�`�b놃d>6=i,K(�!�ą�dZ���^\<�y���V�:�!�W0U0R���,7Q#���⇣N�!�I!5�T�e(!<��� }:!�j5:�"'_ r����ǁX�9!�$
=f�,h�b�?k�DhJ㢞i!�dǹ��dxUD������ʻQ!�� 2]�q�I�969��l��P#28r�"O���G�h�@�5��Ό�uB%D���t�S�f���q�]����j$D�,�NG04����jW/Bɐ(�A�"D�4�t��9�fp3����^EP ��+"D�hHc�U5_d�;"��?]:�0�?D��9�ӵyJ�c��@%"�°&?D���Ե%�<}$k��,�0�a��*D���Ab�X枱��!ш0���'D��ʖȅ������O0u¬�Y�;D�����(P z4#�"4|�~���A9D�� ���=?�!� E
>+NzI�C�5D��Q�k��d����(
4(	�k�g4D���J��&�0�r�b ��as(D�hؠG�F@�0��A� ��Ae%D�,b��B�D!0 
 k2�@e�0D�$a ��0Ƃ ����!��$��g;D�(��6[�z��W'F�z>B�H&":D�x�IԬ���Ҧ�1v�C��9D�̘��m��D�Nޮ@��8D�ૅd�:�b�䯀�n5���׌6D���,W�|�X�k��B�V���2ů4D���voU�-i��AD��&~�\�A�&D�D�T��9m�}��G
F�� D� 0(Fm�� ƨW�d�(� 1D�(����E��@1c�I�x�8�)9D��K2m2n"]�"�u�@	8�8D��Fォdt�$�+���K%�8D����!��v���/��x�t
5D��Q�.B�%�(�r҆ %'�!�D��dAF�P�l�����rgf�Jm!�$N�T����l�$2Z�;�J�=GF!�$�F'x@�4A��a�b�"�I��$!��	2��=@v�� 48�hI:�!��ט2��"�#�Ni敺CȌ��!��ߥ��ՠ�+N�|YF���P�!�$�*S�0P32��pa$,�#n��u�!�ěa��B��y��P�U!k4!�ċ%�>����90�1���-!��Hx$5�`�c>!�$W�f�|0��׮���e��	(!�d�4q(�A�uB��(�P���"j!���?l�I:�Z�,�0��H�!�DH<p9�\j�����&@ϳ`!�DJ8��Y-1c��ӍI�u|a�'b���a�2LX��d�j�
1 �'̀�����S���83I��_Ǻ�`
�'ն�q�����)��g�^Q�q��'}���C�C�`�$hDA�C����'���рN��7t����=Z���'�*�S(�$Na�Æè�j���'\���#M>r�񃳢�39 P;�'�v�{_P���s$@W#`�x��'H��i��3��X�#���&$��'�:�rp/G�dLX�sc����a1�'Uࠁw�h��"���l��'���{ƣÂ�\�2l�=��E��'�㥭O\b�B.�R=��'/�C����h� "B' �0�'���oD;`��9��
�'I~隕Aҙ[X���A�נE>niS
�'
����8���[a�����	�'����F�7�JD�3mė}/h�(�'�Fi�q�D�� �E,	)������ ځ�/ґAt�s�c�Wz�۔"O�b�E@'@�pr5b��ʖ���"O>�wI��\����@��OS"]��"O~��#b��6]�0�H��,�x�� "O9X@f�1��p��&[0D�0����4S���$j���'���X?�r$ŋ�?ӂ��J�Q�6M!`��.=O�8q���?��
Ą`�0"�7��, .�V�6��.k>�P���3A�h�SH��
�X�m%�OB���a�ԺA؄Q`"�s�<�UDH�7\����|?�Aqf��d������'!R� ���?��d�ic.�TLD9���W��h�0F�O��O����O�p��늑8E*��5`�8V�P(A��'�7��O<6����b�� o�'�t���Iı'N�9�I9V]��0ڴ�?����?��'gS��p��?q�4��PID�!e����j��a 蘩5����(1�$��Q	<�֥�'�����X>μI�t�ӌ >
Q�'	�)e�7��/Q�P雐f9�"$QgcA�FoB��;�u�F)���ḧc���>&q)�!P8H,�@�iuH�����?9�O�T�sӆe�O� �؝��E�(4p��O��%�O~� ��8H�$U��h�K��<SW헱osfb����4�?��t�i�~�S��/b���G��:j@1�O����>
�+�C�O>���O0�$�������M3�(+��i�j@	{ ���lG�g��A����� a��ނK���0��O�� Dx���6p¼YD��8դ���h�y�ڸ.ua���MÅz�r�s�b�a��B}��6�TS�$��~a��C���f�c�؃7,��3V|���ȟDyI<�-���g��;�T�I6R��A[,��0�)�矠��NL6� Z��R�p�1�P���r�ҒO�ퟶʓc����2N�jI`l��� ��8@U���*a*� ��?���?	�G͍�?q���?I��:�M���YN�8V�.fp!�f��#������X ��I���Y�'A�}��f��~�P	n��Ȃf�6I�9S�*Vw�yu-��<z7�e��}�?i��Y���l�G�J%h�ꐤU$y��dx0!zǽil2Z��ã	�s�ӺӜO�v]�� �8����Ċr|�5Q	�'�>%B'N���e;`*�6c<L���'�66m����'�J���hb�H�D�O2�'#@x�K���V�(3F���X�0B+T5	��'�b ��ؚ�H�Ɛn|��Oқbnj��'+�t��ٝ3o\��_�a�d Dz'�	Vl���V

vp��۰@]�֝�N\d՛ i^�W��[�L0�$���[`��&������N|��4�5 �E_�3���j��ML���'L�O?��� g��� �ѕ.�ZI�#aE�@иD{���nj��'$��ݢ�+�*w�E ���J����?��3GX� ��r�t!��3(�'���n��`Y�,�������`����V�4��C�+�tZqK�,Ay�@h�I^����P>=���CIX�+b��lĵ���3�����@�A�H��Ɵ"Or�%	�%_��u׾�N]%?�ضe�D�3ͅ�s�=T��<�<7m׈yu��'>�6�O�#~nڈ+���E�&(
�er��c���I� �?��d{"ꁻ�)�?��(��jK%�Q����4�6��`���H�?b�"�r�ʣ~�M��#׾���=	�eT   �   ]   Ĵ���	��Z�Zv)Ċ;R��(3��H�ݴ���qe�H~-�8L,<���i�n�?
.Q�0�đmz(�Ӥ�._6��)�4<�>��' ��0O��@6�ʖ���:"m�&To�pS�Y2j��RߴZBqOR����D^*�MW�[	A�Ʃ+oY�Y��,���V���D 8Qf}I�4$���.�응e�:ל�;R}��c��e�Hu�Ҏ��K$ ����6)<��'���v�Z&(%�OR�2d��v�4�
��ȜJ���ʡ��g��o�$�?i�'Ed���=Q�)-O,��U'J�D��\c�(y�S菳tT,hĭG�WĂ)�O>��M8�zrF�O�mےl�&�,a�fg� M-BA<O��������OH�h2CS"g(�\�-�A��$�r�p�'��IExbkN}�)�?-|���!�T'.��Q�L���W��3F�D� )�����%ߖSjՙ��ʈ.
��J�A�'|ZuDxR���3�|PS�C�����tf6yӨm�}rBK�'�N4䧭<�rME�{�X`�b�,v~�l(O��9��D�<��'}l8�Q�20*i���5g� \A"�V~�'�%Ex��Vߟ�	wA̙D���1!.��8n��X!.&�I�8��x��x����w4����4zxӤ�\.�~R��x�'��(Eyr.ԱtCDI�s�M'�`R���?i$�d}B�8����t��u7:���*eB��t� GOR(�P�H�ƇN�7D,�O�%���\�'}����C]~��t#��� g͌�	4��M>�d�ۈ*6�Q�<�I�)�Xa�(Y�=lT�fЯ�PX��'Nl��@ ��"O��Y�N-W*`���R	Hܩ�D"O��h�f�;P�&�@2�"x�a�3O��x��� K�JQ���ʤl������f���D�4�O�jR'�j�V(�l�P�.��u�	�]�9r��B�T��O:���b�F�44X�(v U����'Q�����3!pĸ��EY�N��I��O��C&��,��l�m
T>��¦��@t�r�lF>]���pH5D��"�/[(j��	���Ĳ���YRL�/O،hVc��9:`<%>c��;��&���į�%!Fb1�-'�O���פ��]i�]k�f�:�%KPN"�í2���B�'�~}i!`�'j[+��I&A�����)��X�KY[���O�q)T�ڱD�� s-�E��-��'aL��⊯\�-3%�>�fix�Ox�Ұ�X�/��If�[>a�    �    R  �  �  &&  x'   Ĵ���	����Z�/C�'ll\�0�|r�'a�	�Dط8��0b�
�<�}#�'�t4��B�h�dt,�:?������i"x�	�-��K����1Bʚ�HH�� Ҕz�J�[�.�0�|)`��u䨉:�Œ�_2Ii�$]�-��s�	��	-�i�V���LX��92��6�x)����sA�)(E&X�9צ��
����q�`˯do���ЂL99}�4y2�E�C����>��(J�"���U�i�����m�<�e���Vk�$�r���3�,���E^�<�Ѝ3?�0���x"���,�]�<�BcQ�P�nЈ�"R�	cT����M�<YDc�r��1��Y�����F�<Q�ձP�҅����*
8�P{6�B�<鲆
(z8���J�%~A�C�N_�<1�!+��|�p!O!gƖkB�F�<��o	�;��B��[;Q�xYq��~�<�և�+}xe薋���b��d�Qf�<�!��.0� �a�=5l���
d�<��"Ι%yMX$(��^W$���|�<I$l[?E~*�l�!Ha�T�C�y4xF~8i�bL�qȂp���y�)�	{O�|���
�txf���J�ym �}Y�*#*��7\�@V$C7�y�M+,:Ѐ�JB�9�0C�gN�y(�q�:�$�M⧄VG!�T'!w���3�X,B���]!�LJ�.h�wD	�6�a�P��(v(!�D4 ���H�o"ʁY��ѻt�!�$!W[V��1΀! 1��F_Z�!��T�Ms�@�/��j���wFòk�!��D��(��&o��B�/E�!��q�%��O�2�&yz�΅�k�!�D��6��<	o�R�(�`�M�<!�ĜRq���Wc&V��K�-<!��yy�����b$�Њ�t/!��H�fؠ���0�����V9!�C�p}܈r�j��Se<���Α�B䉭W����KD��	 �3|pC�"Oh�q[�	 �j�h]j5�փO-�C�I�"�� �S������0��C䉴([4��BH
C��]�2���1˨C�I�3��c0�N�j��q��&����C�ɸ���[2��1-�Q&�̧:�bB�I.t*�]�7+W(8C�[�/Р"�2B�I�r�@�D ���H2���
B�UCL�⋀2:*�b�;|�C�IRU@��m�	8���k��M�BB�	/���ck�u���"D��!:�C�	8W%����o c~�E�D�î�C��
=�x�0�E��-"0�ˆ��7D�fB�	�+���ħ�bm�V�D�y�hB�I;=���+� >�@�1/�4+%XB�	�~0��ԧ�3[i.i�0(��sxB�I,\ ���d�ѵ3!b���S�BB��9�0H��� C'��Bh��)�C�I\���ao� �Ď���C�	;A�d5`���/}����C�(%�C�ɯmh|dZpe��o��0��-�eA�C�	��f����N�h�\�'F�B��C�ɣ;���{LG�s�r�
fσ�l(hB�I�v!��đ$8)F��� �Ju8B�ɣ�dX�g$�6%"��P�S�&Z�C�	��PE�e3}�]�g"ݯ~��C�I>�a��"�1zr6���"X3ZB�I!^0���"#�-<����DX�L�B䉛jwL��JݳM]�X%��`8nC�)� RL�6g\�F�
��f�%Z�"OmQ�2����w	I.80��"O����,���"��c�N�3"O�U��M�B��L�sȞ�M_r���"O��V�>n�A�l&X]+q"Ox In�>�j���	��v�lA@"O��Ct��C�����4E�f�+E"O��1�ED/Cb4�����`)1�"O(� ��bR�@��0���1"O��1BոL�|<"<H�Hq� "O�k��&S<EQ��-���%"O� AqВZ�RP�%����S�"O���cLa6���\Ȉc"OJ0� &Q�z��@I��[�_|��"O��V���:C�t��GB�U�p�i�"Oͨ�k�7���s'��1�U[a"Ov�+v-N3�j@��e�[ߚl� "OZ�b/2�tC1�M�dȞE�r"O8��O�#3�)YE�R5`|�e"Op�ʖA���8�f	�}���"OB�xT�L�P�a��7�%!�"O�8ش��)��t��닦,c�}�3"O�)��M͜�� ��JկZ]�3"O(���	�*�\XtI�xJx��s"O�Y[&�K�AT%���E����"O�-��-Q0 ���K@Kۨ\{XS�"ON9�F�'Tࢯʿ;Q$��"O|Uc؋e$�r� � V��}��"OHp�)��.�a�
�%O�� "OH���DG
�B4�q�L?D�<�*�"OJ���
.q�u
�9�>�s"O�K�%\,NHw	ή8����"O6�˗�SfT����/
��h��"OR5�A,!L2��OS1s��3D"O>q�&I�D2��bNح)���%"O��F��1&ʄ�#��t�#q"OX�����IZP�����3�X��"O^�U��ZrΔ��D���"OL�auGH�|�P+�Ů���"O
���Z3R����鑘b%Ъ�"O���*��? �	�hcܬ��"O�{U�;ø$�ceH�e.���"O�)��ٵj�����Q3'V�@�6"O��Ң$B�O��X�j�ܑ�S"O�Ds���4��R�hN�C��D�G"O��U�O
.1���SD�2��"O�$�R�?OH$q6/ҹ~0H0��"O"�SGF\=RY�#�A&�;�"O,hRe��9Lv�]�%�������"O\�s�M�W��	1��)�BP:'"O
y��D��-$�S�0e��Xxc"O��"�'I�pZ~=2�N�:�6(�e"O�1�7Y�i�PO��85����"O�)��͂&�ikw͕9#�2	�r"O���@�R�������'�,�i�"O8ɱa�٣g��U(sA@�t��e��"O2��SƐ(/9�]ЕG��I� 4�"O ��5������&K�h��\�v"OdiD��"y:�3�>*�"O\�K1�H�]
���
:<�P �"O��X��3�f!CvkFq�d[�"OD������RA^��ֈ$�"O������B���sf�G䨚�"O���Q�Y�8�
�{`�϶X1��ڀ"O� <�G�S/N��0��3M�,�R"O�T%*��x�V!z���|��"O�$r�)��=�l�j���
0�2L�A"O8���I�hV��  ���0�.�c"OT9rn��.�{h��e����"Oe�&o�$t*8Y1�9b��"�"Ot���6���b���bVb�XG*Of���̌����h�H��m����'9:ٚ���-�T� ���P���'�hiC�����K�^0�	 �'�>�bH��^�։8`���R�v=��'��5C���t� �:�ڶi�'��@feC,Sf�P���6F� ԋ�'�t�jb凌0��=Yu��Ky��
�'�pB����<4�$	�,O�Y �'P��c�a�7u�,��ۋ
!F��'Z.@3拌5gf%xg/ܟ h1��'�}y�)Z�=$!r�E�A�4�p�'��xx��o�& ���(w���0	�'ђ]yA`�)"N��"���Z�Ν
�'Q�������!��O�_�* ��'����a&N�{���ѷBR�<�'�@�0�c��,#PQ�4,̋L�x=�'�(J ̊�.�@[�`��~X�`	�'�d=`2��R	�mkƃ��w�+�'��� 針ϊ��1�OOTC�'�6�pED[�.�bp�ƌ�X2]�
�'� Yi�%;
*��E�/_k���'�hu�Ǭ	!f��,��a�G��\�
�'Z�T��x���U��͉�'H��#����xИ$�U_	L� �'�z J�*�&j7�ˤ@�6W��;	�' 
u�E��& ����"Ҍ]	z-��'TDQ{�!��_ H��9b�8�'�Xbc	4qw����!�Ϩ��'� �CmK�o�`��g����A��'��)(Eg?z��-�!˻5��mQ�'�<��Gˋ�[�H`��З7'�t�	�'��Hr��33Z�J�a�>#���P
�'@|	H�i2yN�@b@��1�	
�'�B��e�{�vlx������'�a�v!�+�Is�̝�Y
�'��djG� }��Y��K��3�'�v)�!i� 0��́r��$t��	�'L2���B��(�`'� � �"�'ir@�*M<nh��+Q��F` �'�nL�A')���ĉH?����'�d�`�"˘?+�� �h��<���
�'��q0��Ǣ\f���7���3Ϭ`�
�'�f�[���(U��`����#�$[
�'(̪�E�.\ԡ�1
L���j�'~E�s(*�ԋ���O�f���'��yp N�%f�ơ8$�ͧo�`"�'�49�i_���E䋘�8)����']�u{�l� �*�ɠ�3>1��'c4 v��@�T�JC�:�X�B�'� ��K�/��)�s�*9�\�	�'�$�
E`��1�tAYC��(t�	�'�0�j�D#H�<�ӌ/)��tY	�'4�C,O�=�<�g+׊5/���'4)ˁ��,։H��5�`���'X�4���X
G���iB*�o����'>��r�֊.���u����5!�'�A�(ON����NJˤ�+��� ��H��"4	�	۸rb��t"O9iE^�U<Mp֯ϲ=��� `"O�\�v ��0��E�3��\�"80�"OVI�
[�8p6MYG*�<X���"O�a#�+�o�H���F��Q"O+M��l4́1fO��{��W��!���:B���H�"A�ls��ޮ�!��T��*1�	D(y�(e�!���7 ������ß"c(���ʝ�;�L|�Z�����	�U���A0f��M���z�AS5}߈C�ɨ_��y��$��諤�;GO�B�I`�l�s@�"i��C��B�Ɉc]NL	�Y<,p>��B͍!_ B�I�"(����;�J�*ׯʈt��C�I�'q0҇KL�k�Dl�%���7%�C�ɘa6x(f-T��!I�R�JTB�	�no����N<J_ar�D��$)�C�I�~��D��A�$9X�H�3:�(C䉛62l�����:Qs���2A]t8C��
�QČ�uH�m�����4C�ɰ4,�9��/�}�DS��8HC�I:s*�$sB��}��M��	۬<XB��	) l�
�ϗ <TԽʁ�ܝ�\C�ɰw�,02��"M�dq-�#qC�I%A�4��2��=���a��U�[l2C�	kS�"ң?D�9�%�&V�C��#W�
e�aS=)R`�	`�`,(C��
����c�@9H7�1��+�L��B�	�7�V4��KD%���₢͇*��B��pT\���7bJIR5Ν,U��B�ɃG��8�3�WvP�ȳǫ�u�ZC��C�va�pIW6IfX�Y��G���B�ɯ�
���N�:J2&Ѐo�r\�B�I�Y�d����<#d��$�8D�\C䉾7ܴLRG�§:MrӧN�q)^C�I�>e �b,ؘld���a9U�B�I1>�,��<��T�eFL��~B�	��ؘd��l����i˅�xB�ɯwc``BƊ�9j�p�� ��>��C�2do�X�B���d4�u�˙nK*B��#Q��E�E�V�A)<*��\�g�(B䉁R��� iؿ6�+fě4B�B�$\�� ���҃B����M3�C�	L�f�2v!˙{+*����6{&�C��'^������U>Č:a�ȵ{
�C�ɹy`Jpɒ��	d׆��0��2x�C�2w@v�CƬ�-�\�+�f��D��C�0b��a��ϑ4���`�	y/�C��h��b�A9`���;ׂ_&"�LB�ɖ`���p��^33<xu㥍><�&B�	��Eb�J.z�H��h	�y��C�)2�H��L�Go�Q��JC
M�C��<C����E��N ���l��C�	�\<N��#�G�9�n�!���[��C��2w@L\9p'�!&n:�t@�t�C�ɸ�0���H� �5�h ��"O�1i��$a1�%��N#���w"O��။�=�;�N�dnI��"O4��1cM�{jY;��@�~4�[�"O����+U2�>Ds�,1�(�D"O�,��d,
� �LU�e�h��"Or�X7��'�Th�����Ф�e"O��
��ݫ*|�!�*_�{p��"OV���mځ-(Ah���fĭ9�"O� ��Au��!pe�r�#VmC�m�"O��B&D��qQd#)�졐P"O>�&���T�
	�b^t��E	�"O�������l��YG�&���"Ovѓ1IZ�~�B���<���"Or\�Ԉ��Q8��Ǌ!;�"�Ѓ"OL��"A��^�|���}�̴��"O�(��*ٵ5Ȳ]���="1�5"O���#Ip�Q2��E�1�"O�Yk�d��CtCƣ�tzd"O�B���:�d��vǏ��~�"O^�h��!�0�r�EQA�|ZT"O�e�b�Z�E�X�7ś�0�v�;�"O���קÇ ���c4��3	nd�H2"OA���D:]�:�+�dC�WevВ�"O��鐀љS�&�1vAD�j>pd�w"O�Ѱ7O����V�X#���%"O�|�$j�{[`��$��K�80�'"O��c4&ǆuw��'B� j����"ON=�/B�H�ോb� M�1[g"Or�
e���ޕzf���5�
ŨT"O���g ���}�a��6���[�"OB�Z>]����ɋo&lA5"O��2�.ɥ"��E�'��8&�H"O
�O�!|1�$���5W�8S�"O���皅t��p!	K�����"O�(���L}����+D��}h�"Oj`"��
�4YR�VO�"J��"OF]�f'J�~{���Q��-j��"O �#$jJ�& �1t,D�o_��(�"O�$��Z� �:�+��$<:�S"O��Z��7"M �2�X����"O�0rfhR;j��T FfE,�� pt"O<Ձq�٣<a��Җe��|��)8�"O�Q`i��~�˳N�M��E��"O�X��]!j�z�ʲg�$���"O�RQ���:x@�&旯Mΐ�%"Oh83���u���@��1r�b�+�"OBU�&e	�Wr�c5��rߊ%�d"O�[V%�	�00���NΞQ�"O�Ѳ3o[a�D��?mZ�*f"O$�V��/?j�A5BO�gNr�a�"O�Uk�e�xz��O�6C�I#�"O�����״��狊�ba)�q"O�����r8�r��5X����"O����Ώ�*dX�RIƀ@T��`1"O@R�+cq~Sw�֨_>�i�"O�ɘ D	T@��� ̯Tŀ�		�'�J8�Fo_;iQ��HS
�b9�'A*���+�
Z*�S� ��>�+�'�:�u�
~j���rg��	ޤ�'�"�b��$KU,t@��M3���'��8�H��dK��Q1�^~
@��'�hh��Ȃ���yc�ȶ�nL��'�(���8�ԅkU��x���K�'�P8��
LAk���.��h��`!�'��j��^+q����dgN^�4�8�'`�A���{��e񠝉P��h�'=b����b��%
Q�]�LRFD��'���Z&�@G(TK���G� �
�'�|�����<�8� #�P�r���'���5� [�p�oQ
	?Ҩ��'��iD�������E��t��'���hAe�0{A�]�@!��s�"O� ��it�̮w�X#��U�i���p'"O<���F]�h�H����E�)�
#�"O�H2�� &�~ŃW%I�i��8��"Oּ�Q~AZ��A]��M{�"O2`����;�e���<?v&��"Oq@
,0�H���9���r#"Op���h�R��%͜A�X�4"O�bdm��.�n :��¥w|N	sa"Oȅ����~8ȡA1��q�A��"O��S�R�@Ъ�����! X��I�"O�u� �0f�Z=�ꗆe�
pb"O���G&ɶc;���J��t��<��"O�Q�ggd\��(ң=�zm�"OL1���>V���Є�D�bΦpa"O�lS�m��?����W�`�
��"OPy��7	r,P���"�xʆ"O`�������X�=��Y��"OT�ڥ"�*\xi�� g{�,+c"OP�Pq�C�F.6�Z'��^���i'"O�����<O��Ex&�Z�Cy(U˅"O������z��鳒�!<O`�Q"ON���O'Fp����Ȥ[6�-XP"OJ0ˁb�>(��ظE)��T��U��"O�Ȁ�+��*�*%ZI��w���R"O�	
���R��D������c�"O���!ڸ��q*�ǋ�`����"O�䂐�@z�܌���K#����"O0��"��(Ј�j0-º� T"Obh�r�.+�0C����,E�̹q"O�S���|ء�&�$=�}X "O��R�?��[a`��/:� �"O<�;� �=��4�q�_�&��"O�XǤT�t�\A9E�ǒy�혰"O���N� /�0IA%G�u�Yv"O*c�&�t���r�B�T	� �"Oe��!�$9t��f�_�"�|���"OR`rv#LHH�I�i�4B�pLQu"Oڽ���� ^��E	�~�p��"O��AG
�>�>d��g��� �"OB����[�P��d� fU �=�"ONI,,��"Q�**a�*[�!�d�7:�d�V�Q�~�6����T�D�!�Z�A�ܵ��m�	E�bO��!�d��l2��#+�2 :�`��� �!���46(���J&P�y����	W�!��P�o�vMZ�B�|��1���!�C>^�X���{��=��얖o�!�ă�<ۼ�2f���I0=�JD�e!���(A�^� 2�Z�F�l�K��A��!��;wA�\�ש,H�� b�@5!�ϓ(����m�09�P`˽q!�D@�Gl���]�O��`g�1m�!���r5a%+°L{��1�Ơz�!�D
�;@X���N,�[���Q!�$O��$����b�ڠGX�,a!�f� ��X�~_�mA&@�$!�D���l5�#�JW���q���>!��/zV��I��mSԂլ��u!��^�rh����=q��sDMZ�Z�!��5Rz"@�����6DJ�Z
&�!�Ԅ8j  �d'�4D���F�!�$];��!4M�p���Sc�V$G�!����5A&O�R)>=q0$�!�d�6tF�cB�;r�Yc��j!�� �$c D�u�ʌ@�R�5/f�s"ObP�����C"��:P���*�0�`�"O�9�J��:�H�;��&U�
5�P"O���^XI�����9��"O��X&�֕F]�Dm��`=�"O�ŲEK�6=a~ɲ���!J�{�"O4\ɒ��-+V!��%g�#"O�%c�Òr di�Hج<|��"O�� �鄌uܘ�'��O�|�"O�t�/�R<p8���9�@��"O��QV�D�*>�h���"����"O�|Cq
�1�t��$i	(P�zM�2"O��Ы��)�q�Gǉ�SbF��"OB���  �   j   Ĵ���	��Z�RV)Ǒ7>��(3��H��R�
O�ظ2a$?����H�49a��i��I��i� ]�=����V`�6̀��9X�4Z���a�'[�V��p�4�I�8QP�Z�d��V}@����2Sd#<G�5x�67�]�|mN![g
��{� < gÌ,%���`8����2��L�OUrQ��_�qJ��'h�As&N���3�f�p4�+��5��L�?{�L%�z#
1;w�Z�.���ԟ6��6D�	2K�*ְ���qn<!(��C�+R!" �O�� �%�W`6�h�X�����<���� D�>b x�֍_�Ԓ�-[�2$R��'׮���d	@�'���'�)��N�6"� mԈv,�4rhe��i��I"5��H�/X)c7�!B-�2N$K' 8�O���Ď#��� [��e�@X1$s�����L)tg�H#<��6�Iƒ�l�D�<\:��iМ�B��i�qDx�k�L�'�t�dW5@eĸ3ڳ<=��IY��'pz�Ex�p~�JÝi!��p�A�Q4��[5�ի��$�'�O������,-d�FB��L�2�H��خ7�4Ex���f�'D�!�I#e����0fZ ���C�6h$�b�( G�I�'{0�PrNЀv�(0pC�D�441�'}HDx���I8[���fKG?�d��fc��e���T�ۚ,>� �%o��Y+ߴRk�|CCJG�'t��*����u��ߢ&XTx�@�ڈI�DX۔
�^qORl���[
����X��ǈa� �:Ή�7�P��%X6�q'����(O<U��ҳf����Ϩ(2���"O,���  ��]�\	.#�p�A*��Ɇ4`�(�b�V����hR��LmJ��B�&��G=�¡:Wid�E�CF"t�p�җ#�3u�	���M��$@# �<��h
93Q�����-A"Kc�\�"�O��0«?D�0�k�%k�r��"T�]v�ʀL�<��'�B�0gTd
̀1႕19J"ܮj�FDB�'m���@��|ɠmҋV&X��דj�2i��)b��;����F�H��3?e{�N��2W��# b�Gٹ_�<A��cy���3�j��M(����$���	�� �=��$ ̐P��gR!:��I""�L|�#h�29�B䕴f�y��_�C:9��#���?Q�HA*1��J�\?��,p�e�����4����ݲ�(O�t��S��,
�8    �    R  �  �  &&  x'   Ĵ���	����Z�/C�'ll\�0�|r�'a�	�Dط8��0b�
�<�}#�'�t4��B�h�dt,�:?������i"x�	�-��K����1Bʚ�HH�� Ҕz�J�[�.�0�|)`��u䨉:�Œ�_2Ii�$]�-��s�	��	-�i�V���LX��92��6�x)����sA�)(E&X�9צ��
����q�`˯do���ЂL99}�4y2�E�C����>��(J�"���U�i�����m�<�e���Vk�$�r���3�,���E^�<�Ѝ3?�0���x"���,�]�<�BcQ�P�nЈ�"R�	cT����M�<YDc�r��1��Y�����F�<Q�ձP�҅����*
8�P{6�B�<鲆
(z8���J�%~A�C�N_�<1�!+��|�p!O!gƖkB�F�<��o	�;��B��[;Q�xYq��~�<�և�+}xe薋���b��d�Qf�<�!��.0� �a�=5l���
d�<��"Ι%yMX$(��^W$���|�<I$l[?E~*�l�!Ha�T�C�y4xF~8i�bL�qȂp���y�)�	{O�|���
�txf���J�ym �}Y�*#*��7\�@V$C7�y�M+,:Ѐ�JB�9�0C�gN�y(�q�:�$�M⧄VG!�T'!w���3�X,B���]!�LJ�.h�wD	�6�a�P��(v(!�D4 ���H�o"ʁY��ѻt�!�$!W[V��1΀! 1��F_Z�!��T�Ms�@�/��j���wFòk�!��D��(��&o��B�/E�!��q�%��O�2�&yz�΅�k�!�D��6��<	o�R�(�`�M�<!�ĜRq���Wc&V��K�-<!��yy�����b$�Њ�t/!��H�fؠ���0�����V9!�C�p}܈r�j��Se<���Α�B䉭W����KD��	 �3|pC�"Oh�q[�	 �j�h]j5�փO-�C�I�"�� �S������0��C䉴([4��BH
C��]�2���1˨C�I�3��c0�N�j��q��&����C�ɸ���[2��1-�Q&�̧:�bB�I.t*�]�7+W(8C�[�/Р"�2B�I�r�@�D ���H2���
B�UCL�⋀2:*�b�;|�C�IRU@��m�	8���k��M�BB�	/���ck�u���"D��!:�C�	8W%����o c~�E�D�î�C��
=�x�0�E��-"0�ˆ��7D�fB�	�+���ħ�bm�V�D�y�hB�I;=���+� >�@�1/�4+%XB�	�~0��ԧ�3[i.i�0(��sxB�I,\ ���d�ѵ3!b���S�BB��9�0H��� C'��Bh��)�C�I\���ao� �Ď���C�	;A�d5`���/}����C�(%�C�ɯmh|dZpe��o��0��-�eA�C�	��f����N�h�\�'F�B��C�ɣ;���{LG�s�r�
fσ�l(hB�I�v!��đ$8)F��� �Ju8B�ɣ�dX�g$�6%"��P�S�&Z�C�	��PE�e3}�]�g"ݯ~��C�I>�a��"�1zr6���"X3ZB�I!^0���"#�-<����DX�L�B䉛jwL��JݳM]�X%��`8nC�)� RL�6g\�F�
��f�%Z�"OmQ�2����w	I.80��"O����,���"��c�N�3"O�U��M�B��L�sȞ�M_r���"O��V�>n�A�l&X]+q"Ox In�>�j���	��v�lA@"O��Ct��C�����4E�f�+E"O��1�ED/Cb4�����`)1�"O(� ��bR�@��0���1"O��1BոL�|<"<H�Hq� "O�k��&S<EQ��-���%"O� AqВZ�RP�%����S�"O���cLa6���\Ȉc"OJ0� &Q�z��@I��[�_|��"O��V���:C�t��GB�U�p�i�"Oͨ�k�7���s'��1�U[a"Ov�+v-N3�j@��e�[ߚl� "OZ�b/2�tC1�M�dȞE�r"O8��O�#3�)YE�R5`|�e"Op�ʖA���8�f	�}���"OB�xT�L�P�a��7�%!�"O�8ش��)��t��닦,c�}�3"O�)��M͜�� ��JկZ]�3"O(���	�*�\XtI�xJx��s"O�Y[&�K�AT%���E����"O�-��-Q0 ���K@Kۨ\{XS�"ON9�F�'Tࢯʿ;Q$��"O|Uc؋e$�r� � V��}��"OHp�)��.�a�
�%O�� "OH���DG
�B4�q�L?D�<�*�"OJ���
.q�u
�9�>�s"O�K�%\,NHw	ή8����"O6�˗�SfT����/
��h��"OR5�A,!L2��OS1s��3D"O>q�&I�D2��bNح)���%"O��F��1&ʄ�#��t�#q"OX�����IZP�����3�X��"O^�U��ZrΔ��D���"OL�auGH�|�P+�Ů���"O
���Z3R����鑘b%Ъ�"O���*��? �	�hcܬ��"O�{U�;ø$�ceH�e.���"O�)��ٵj�����Q3'V�@�6"O��Ң$B�O��X�j�ܑ�S"O�Ds���4��R�hN�C��D�G"O��U�O
.1���SD�2��"O�$�R�?OH$q6/ҹ~0H0��"O"�SGF\=RY�#�A&�;�"O,hRe��9Lv�]�%�������"O\�s�M�W��	1��)�BP:'"O
y��D��-$�S�0e��Xxc"O��"�'I�pZ~=2�N�:�6(�e"O�1�7Y�i�PO��85����"O�)��͂&�ikw͕9#�2	�r"O���@�R�������'�,�i�"O8ɱa�٣g��U(sA@�t��e��"O2��SƐ(/9�]ЕG��I� 4�"O ��5������&K�h��\�v"OdiD��"y:�3�>*�"O\�K1�H�]
���
:<�P �"O��X��3�f!CvkFq�d[�"OD������RA^��ֈ$�"O������B���sf�G䨚�"O���Q�Y�8�
�{`�϶X1��ڀ"O� <�G�S/N��0��3M�,�R"O�T%*��x�V!z���|��"O�$r�)��=�l�j���
0�2L�A"O8���I�hV��  ���0�.�c"OT9rn��.�{h��e����"Oe�&o�$t*8Y1�9b��"�"Ot���6���b���bVb�XG*Of���̌����h�H��m����'9:ٚ���-�T� ���P���'�hiC�����K�^0�	 �'�>�bH��^�։8`���R�v=��'��5C���t� �:�ڶi�'��@feC,Sf�P���6F� ԋ�'�t�jb凌0��=Yu��Ky��
�'�pB����<4�$	�,O�Y �'P��c�a�7u�,��ۋ
!F��'Z.@3拌5gf%xg/ܟ h1��'�}y�)Z�=$!r�E�A�4�p�'��xx��o�& ���(w���0	�'ђ]yA`�)"N��"���Z�Ν
�'Q�������!��O�_�* ��'����a&N�{���ѷBR�<�'�@�0�c��,#PQ�4,̋L�x=�'�(J ̊�.�@[�`��~X�`	�'�d=`2��R	�mkƃ��w�+�'��� 針ϊ��1�OOTC�'�6�pED[�.�bp�ƌ�X2]�
�'� Yi�%;
*��E�/_k���'�hu�Ǭ	!f��,��a�G��\�
�'Z�T��x���U��͉�'H��#����xИ$�U_	L� �'�z J�*�&j7�ˤ@�6W��;	�' 
u�E��& ����"Ҍ]	z-��'TDQ{�!��_ H��9b�8�'�Xbc	4qw����!�Ϩ��'� �CmK�o�`��g����A��'��)(Eg?z��-�!˻5��mQ�'�<��Gˋ�[�H`��З7'�t�	�'��Hr��33Z�J�a�>#���P
�'@|	H�i2yN�@b@��1�	
�'�B��e�{�vlx������'�a�v!�+�Is�̝�Y
�'��djG� }��Y��K��3�'�v)�!i� 0��́r��$t��	�'L2���B��(�`'� � �"�'ir@�*M<nh��+Q��F` �'�nL�A')���ĉH?����'�d�`�"˘?+�� �h��<���
�'��q0��Ǣ\f���7���3Ϭ`�
�'�f�[���(U��`����#�$[
�'(̪�E�.\ԡ�1
L���j�'~E�s(*�ԋ���O�f���'��yp N�%f�ơ8$�ͧo�`"�'�49�i_���E䋘�8)����']�u{�l� �*�ɠ�3>1��'c4 v��@�T�JC�:�X�B�'� ��K�/��)�s�*9�\�	�'�$�
E`��1�tAYC��(t�	�'�0�j�D#H�<�ӌ/)��tY	�'4�C,O�=�<�g+׊5/���'4)ˁ��,։H��5�`���'X�4���X
G���iB*�o����'>��r�֊.���u����5!�'�A�(ON����NJˤ�+��� ��H��"4	�	۸rb��t"O9iE^�U<Mp֯ϲ=��� `"O�\�v ��0��E�3��\�"80�"OVI�
[�8p6MYG*�<X���"O�a#�+�o�H���F��Q"O+M��l4́1fO��{��W��!���:B���H�"A�ls��ޮ�!��T��*1�	D(y�(e�!���7 ������ß"c(���ʝ�;�L|�Z�����	�U���A0f��M���z�AS5}߈C�ɨ_��y��$��諤�;GO�B�I`�l�s@�"i��C��B�Ɉc]NL	�Y<,p>��B͍!_ B�I�"(����;�J�*ׯʈt��C�I�'q0҇KL�k�Dl�%���7%�C�ɘa6x(f-T��!I�R�JTB�	�no����N<J_ar�D��$)�C�I�~��D��A�$9X�H�3:�(C䉛62l�����:Qs���2A]t8C��
�QČ�uH�m�����4C�ɰ4,�9��/�}�DS��8HC�I:s*�$sB��}��M��	۬<XB��	) l�
�ϗ <TԽʁ�ܝ�\C�ɰw�,02��"M�dq-�#qC�I%A�4��2��=���a��U�[l2C�	kS�"ң?D�9�%�&V�C��#W�
e�aS=)R`�	`�`,(C��
����c�@9H7�1��+�L��B�	�7�V4��KD%���₢͇*��B��pT\���7bJIR5Ν,U��B�ɃG��8�3�WvP�ȳǫ�u�ZC��C�va�pIW6IfX�Y��G���B�ɯ�
���N�:J2&Ѐo�r\�B�I�Y�d����<#d��$�8D�\C䉾7ܴLRG�§:MrӧN�q)^C�I�>e �b,ؘld���a9U�B�I1>�,��<��T�eFL��~B�	��ؘd��l����i˅�xB�ɯwc``BƊ�9j�p�� ��>��C�2do�X�B���d4�u�˙nK*B��#Q��E�E�V�A)<*��\�g�(B䉁R��� iؿ6�+fě4B�B�$\�� ���҃B����M3�C�	L�f�2v!˙{+*����6{&�C��'^������U>Č:a�ȵ{
�C�ɹy`Jpɒ��	d׆��0��2x�C�2w@v�CƬ�-�\�+�f��D��C�0b��a��ϑ4���`�	y/�C��h��b�A9`���;ׂ_&"�LB�ɖ`���p��^33<xu㥍><�&B�	��Eb�J.z�H��h	�y��C�)2�H��L�Go�Q��JC
M�C��<C����E��N ���l��C�	�\<N��#�G�9�n�!���[��C��2w@L\9p'�!&n:�t@�t�C�ɸ�0���H� �5�h ��"O�1i��$a1�%��N#���w"O��။�=�;�N�dnI��"O4��1cM�{jY;��@�~4�[�"O����+U2�>Ds�,1�(�D"O�,��d,
� �LU�e�h��"Or�X7��'�Th�����Ф�e"O��
��ݫ*|�!�*_�{p��"OV���mځ-(Ah���fĭ9�"O� ��Au��!pe�r�#VmC�m�"O��B&D��qQd#)�졐P"O>�&���T�
	�b^t��E	�"O�������l��YG�&���"Ovѓ1IZ�~�B���<���"Or\�Ԉ��Q8��Ǌ!;�"�Ѓ"OL��"A��^�|���}�̴��"O�(��*ٵ5Ȳ]���="1�5"O���#Ip�Q2��E�1�"O�Yk�d��CtCƣ�tzd"O�B���:�d��vǏ��~�"O^�h��!�0�r�EQA�|ZT"O�e�b�Z�E�X�7ś�0�v�;�"O���קÇ ���c4��3	nd�H2"OA���D:]�:�+�dC�WevВ�"O��鐀љS�&�1vAD�j>pd�w"O�Ѱ7O����V�X#���%"O�|�$j�{[`��$��K�80�'"O��c4&ǆuw��'B� j����"ON=�/B�H�ോb� M�1[g"Or�
e���ޕzf���5�
ŨT"O���g ���}�a��6���[�"OB�Z>]����ɋo&lA5"O��2�.ɥ"��E�'��8&�H"O
�O�!|1�$���5W�8S�"O���皅t��p!	K�����"O�(���L}����+D��}h�"Oj`"��
�4YR�VO�"J��"OF]�f'J�~{���Q��-j��"O �#$jJ�& �1t,D�o_��(�"O�$��Z� �:�+��$<:�S"O��Z��7"M �2�X����"O�0rfhR;j��T FfE,�� pt"O<Ձq�٣<a��Җe��|��)8�"O�Q`i��~�˳N�M��E��"O�X��]!j�z�ʲg�$���"O�RQ���:x@�&旯Mΐ�%"Oh83���u���@��1r�b�+�"OBU�&e	�Wr�c5��rߊ%�d"O�[V%�	�00���NΞQ�"O�Ѳ3o[a�D��?mZ�*f"O$�V��/?j�A5BO�gNr�a�"O�Uk�e�xz��O�6C�I#�"O�����״��狊�ba)�q"O�����r8�r��5X����"O����Ώ�*dX�RIƀ@T��`1"O@R�+cq~Sw�֨_>�i�"O�ɘ D	T@��� ̯Tŀ�		�'�J8�Fo_;iQ��HS
�b9�'A*���+�
Z*�S� ��>�+�'�:�u�
~j���rg��	ޤ�'�"�b��$KU,t@��M3���'��8�H��dK��Q1�^~
@��'�hh��Ȃ���yc�ȶ�nL��'�(���8�ԅkU��x���K�'�P8��
LAk���.��h��`!�'��j��^+q����dgN^�4�8�'`�A���{��e񠝉P��h�'=b����b��%
Q�]�LRFD��'���Z&�@G(TK���G� �
�'�|�����<�8� #�P�r���'���5� [�p�oQ
	?Ҩ��'��iD�������E��t��'���hAe�0{A�]�@!��s�"O� ��it�̮w�X#��U�i���p'"O<���F]�h�H����E�)�
#�"O�H2�� &�~ŃW%I�i��8��"Oּ�Q~AZ��A]��M{�"O2`����;�e���<?v&��"Oq@
,0�H���9���r#"Op���h�R��%͜A�X�4"O�bdm��.�n :��¥w|N	sa"Oȅ����~8ȡA1��q�A��"O��S�R�@Ъ�����! X��I�"O�u� �0f�Z=�ꗆe�
pb"O���G&ɶc;���J��t��<��"O�Q�ggd\��(ң=�zm�"OL1���>V���Є�D�bΦpa"O�lS�m��?����W�`�
��"OPy��7	r,P���"�xʆ"O`�������X�=��Y��"OT�ڥ"�*\xi�� g{�,+c"OP�Pq�C�F.6�Z'��^���i'"O�����<O��Ex&�Z�Cy(U˅"O������z��鳒�!<O`�Q"ON���O'Fp����Ȥ[6�-XP"OJ0ˁb�>(��ظE)��T��U��"O�Ȁ�+��*�*%ZI��w���R"O�	
���R��D������c�"O���!ڸ��q*�ǋ�`����"O�䂐�@z�܌���K#����"O0��"��(Ј�j0-º� T"Obh�r�.+�0C����,E�̹q"O�S���|ء�&�$=�}X "O��R�?��[a`��/:� �"O<�;� �=��4�q�_�&��"O�XǤT�t�\A9E�ǒy�혰"O���N� /�0IA%G�u�Yv"O*c�&�t���r�B�T	� �"Oe��!�$9t��f�_�"�|���"OR`rv#LHH�I�i�4B�pLQu"Oڽ���� ^��E	�~�p��"O��AG
�>�>d��g��� �"OB����[�P��d� fU �=�"ONI,,��"Q�**a�*[�!�d�7:�d�V�Q�~�6����T�D�!�Z�A�ܵ��m�	E�bO��!�d��l2��#+�2 :�`��� �!���46(���J&P�y����	W�!��P�o�vMZ�B�|��1���!�C>^�X���{��=��얖o�!�ă�<ۼ�2f���I0=�JD�e!���(A�^� 2�Z�F�l�K��A��!��;wA�\�ש,H�� b�@5!�ϓ(����m�09�P`˽q!�D@�Gl���]�O��`g�1m�!���r5a%+°L{��1�Ơz�!�D
�;@X���N,�[���Q!�$O��$����b�ڠGX�,a!�f� ��X�~_�mA&@�$!�D���l5�#�JW���q���>!��/zV��I��mSԂլ��u!��^�rh����=q��sDMZ�Z�!��5Rz"@�����6DJ�Z
&�!�Ԅ8j  �d'�4D���F�!�$];��!4M�p���Sc�V$G�!����5A&O�R)>=q0$�!�d�6tF�cB�;r�Yc��j!�� �$c D�u�ʌ@�R�5/f�s"ObP�����C"��:P���*�0�`�"O�9�J��:�H�;��&U�
5�P"O���^XI�����9��"O��X&�֕F]�Dm��`=�"O�ŲEK�6=a~ɲ���!J�{�"O4\ɒ��-+V!��%g�#"O�%c�Òr di�Hج<|��"O�� �鄌uܘ�'��O�|�"O�t�/�R<p8���9�@��"O��QV�D�*>�h���"����"O�|Cq
�1�t��$i	(P�zM�2"O��Ы��)�q�Gǉ�SbF��"OB���  �   \   Ĵ���	��Z�v�G�4P��(3��H��R�
O�ظ2a$?�K&����4`��b�wa��2�� l�B��"#^
�7��Ԧ={�4C�2���:�'��&��(� ��8 �� �L6xT��B��v�`Od��� 0�O��_=	`�@�NC�^�p��Fꋈ	�,ё�\Cy®A�����tgI�����)\j�)�6�����W�8=F�k�΀*d�`g�,}�z1s���<��$។A�T)O`��D�ֆ ��T�ˬS���3Ҫ]!x3��� �x2��w�b�����$��'j���'�n�"�<bΪ!��EBdiBL��P��r�O-P�Q�(��|b�ҦL�x�@�Ѳ.�`�����yOOX�'f�FxB�7� \�%BQV4�p��7��#<��-�a�"� �,i���6H"rlH]��d�O�mh��?�'+���f^.D���������Rݴk^,#<	u-4�j�P���mU�}�ƜJW��Yg��q�Q�F��#<��h!?� �`�J՚��>\�����`�Gy�dVD�'Z�0�?�R-��	�sݏ���Ќ�Qլ#<�0J%-��d}50!X��[��3�ߌ�1O�#��D�!��Y��т&����h�@�>
��@��6Ŋ#<y�F'�I��
^9���;� JDb�S��'���ӯO"�y"�(_�1�|aa���y�×�#z��0c��;*���Dj����/P��r�|⍗> �@J<Q�*.rcJ%
�G �?H��MW�3���rTf�e�	h1r�C��4�Ie꼼��U9%��Řu�Ȝ�c��XB��;��  �$��U�<��C>A�qt�V5��|hG�g�<�@cE�0a��+z�8w+�K�<qTaU�D��p�lФ_z�����G�<a�'־P�b-�T�P>�(�@�G�<a 
(@͒�z .��?
��1�j�n�<��&=lH i�bI9B�!���n�<Ir�ƛ4�̈@���!p�!@i�<���Ÿi]L�#J�P}�����b�<IRB��"�!��	�Ĩ�wD�^�<���8p 4�J�u�N�Cv��Z�<� E�d�Ҏ��!`�� y��RT"O�p[ŧ�޼A�4�@m�^\��"OX��H �2!z�� � z@dxҔ"OF$�U�ܳ3�D���h�7|�jp"O�;� \\�01�G�	���9"O�	)����,-�p����R��A"O���f$�>Bx�)���	��"O�   �  o  �  �  f%  .  K4  �:  �@  G  WM  �S  �Y  `  _f  �l  �r  (y  i  ��  ��  3�  v�  ��  ��  x�  �  �  �  ��  +�  ��  ��  4�  (�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;����i`9"�ˁl�$@��- G��D��O��2�	!0L�Qd�*��PZg"OJ�R������qE����Li�"O@ӥg$x�|���ֱE{�Q�"O��"W����i��ۇI<���"O4)遪@7��P�����z:�!Y"O6�#�`��U�|����%(@"O��J�΅-����		���	շi�hC�I�(���Q7n׭A)�� ���G22B�	�{n@ 8%�@��j�;(��!@�C�	�/���#�"[���@(K�c�E{��� &a����k)�
Da��>�~���"O����<A)
H�B�%`��i�w"O̕(K*$r�"�d̩�XС�"O� �fn�-V�&�
C$M&0��RT"O���T�'7_�����߇ke:%��"O\6�&un���'��V��
��6D��xr�@�I�H�j�O
<��x��"4�	}���Oi�s��Ki����Q�7
XJ�'��|A���{JT���5�
�b�'^d	�u�Y<��k��}e>e[
�'*j�� ��,3`��{�[u�m�ش�Px�E7Q�I�T�[�\���)ȫ��=���|�!�-%Z�xf�@�N��P�d���y�E�0P�ܐ��K(L���;R����'cў�Oz4�c�Z>��H
�B�Pu����'���e	ݬG�.� ��>P���'� ؐe
T	v� p��_�R;�'��<��ǔ&�v*�)T�AL���#��;"� JC@�X��L9,0�@��"O�u��"FKT�D� �ԧ}�h$""O�h"'�;Hs�Sdd��op���'Vў"~��&L(
m��nS;#g���¡X��y�W�z�B)�֡ڞ$�.�������yH�jT��ߑ1�%R���0�yFR�5X��]�$��,���y�)�6{���Fj\9N9bT���X6�yb��@f�\�Z�RC�߀�y"��KN<�P�O��+J� ����0<Q����)+TX�i�)�d7�����Q�]�!�E�8���P�	�<F٢6쓃$֢=E��'-����@,S�b��7��`H$z�'���/�r� #TfΞfE8yK��?	� ��3��.BD3v�/�>����H�MY�قG�1c?zib�e�8ʒB�$q�zA�''�m�L�?J�|��O�"~J���/�  �@�ӫ�"J�I^I�<	e�)�8D�A���MM\�	PdC�'��yr,G������C&�Zr�E��y2]%B�F��S.˚<�`�Z⡐�y�����������"1��أQ� >�O	�'NQ>9�0װk��18�)+u~mɧ!$D�����p#ȰR(�<=ެ��Se�hO�Sb�)�Ma�
R	��Ԡ�LK2�U��nNZxB��nՖ` ��5�hd��O*]
R�Ӵ �ia�F�GbJq���D���,i�i��9+��PC����!�M1Yl�)rfA�L�L=�H]�!��	4��a��,ۊ_C�ecwf�<{o!��B��j�S�ȧf#�p�$F݌5X�^�h�<E��4O���"$%U8���Ýzsb��ȓ]�~�bh��J��1�SZ��}�ȓ
V���`ǔ1J	9e�O.�8e��I�
�v�R��Tي@M҄�����ޔ�y��=R1��Q�>�<$��8�y�n�e�Js�"G��h 1aU"�y�d���Y��)9&�]��2�y��� ��U$�.;�虹#A��yˇK7`˱��_�p����yRF�&s�L�X���N��y�6eǍ�yD��{˒��F��� z|:����y"A�;p!��`�VΌ���'�۰<���̵~����A3?��!
�����!�Dә~�X���L�.�xIyVQ�c�!��\���8ׁ �<�.D�C˅�z!�� �B���ndt� "G�T�tR�"O�LB &t��]ZP P/O#N[�"OA�Gx�����l��I,�a��"Ol�����-! �@��I&3t���"Oz��e�(o�2E��gH��1�"O5�1�+>ꂬ��L��_�e��"O`��5��#J�)�3��(�֩�"O�=�s!�c^t� S)�q�Dɂ"O����v�n�Kc�������"O1:3���,8�u�@�S1�ّ�"O�xjW���4�<��1ę
*����'���8���\y��`,A�i� h��3D���i1)��K׋Jd��TR"G/�nӺ#<�}�PB�d��Ђ҅�F��a]@�<��k`����q�]x�t����Q�'��yrj9
�ہ�ĕI��ڥ%�(�yں�v]+P�J vM�8����y¨�Q���
�>k_ ����ybD٬Z���@gG1cpuZ�ɔ�y�m����J��@6k�`:'˟)�y򣀿��U�F�ZmyrP�L��yBf��=~���cV-c�4-�F�&�y"�m�11p �)^[.�ň϶�y��K/�9Jpd�JЬ��)��yB./M��}���2F���# ��y-�*�	��7�������y���8E�Er3���'����D��yB��k�<��w�"��ӬC4�y"��/7X�RD�j�J-�r��y�7U��)&̒?s��2L^-�yR�H��U���X�W�$�h#S��yR"�D6�E�&~��E���y�L��14��2咿"7D���
�7�y"GE�� �#��.J�Q�K��yrN�9Y��:ebR���U8!��yRE�]�}Y�!~J� :����yr��=	NI�u�D�!�8ʗ��4�yHI6�zb!�	���Y ��7�yR��r�V�����
>��H���y2��" ��ܒ��ԛ"p�����yR�
!J�f�Y��	�\IҊ�0�y���f��2L�
㔍k��A��y�F�:sx��+�����siC �yҊؑ��M�2�� r�X �m�yb�5a�e���X�.��*��y���q�| :�腼9ْ� ��yBEϺI��Ȉ&�֗8<�@�F<�y���(H#�X�z?(�zP�Z�y��(E�0%V�K�C.�21ې�yb�D�Q&�۷��8J&u���)�y�x�X��膛9����
�ybE�f���%�h΀����y�k?i�̺Qώ>=������yR/
g��@z�c�!e�(�]1� B��.O������tm��җ+"RB�I�~5�wHP�Y ��V�V�NUB�ɁRRͻ׆�"*�T&¿U�C�ɳ(��LPU�S��Y�_J��C�	�tx�QB̗A��c3bX/)��C�I*aC�]��Fߒs��5Hv}FB䉀5�����i~k�ꔟqQjB��K%{�`�>m墵�B`_(/ݤB���A`�.O��F�
���3�xB�I%�!+��X�Fi<���Έ,,$(C�)� J�c�O;}n-�$�N8E��i!"O��z@��t�N'@K�h��q ""O�*3쓳1�	�C)�2�@�9�"O6tA�͕�)�A�'>�=��"O �0"�Mb�%��8[y���'%�'���'$��'e��'s��')ґ��  Tz��# ��vX�4'�'��'���'w��'e��'^��'*���)߁9]N�����<V�QW�'���'���'o��'c��'"�'�|�Y�Η0{���6
��j � ��'���e�i%��'�R�'���'f��?t�X�(s,N9j2S�@���'���'��'b�'���'�b�'݀<
�^�Aڰ����Ɓt�"�b��'cr�'CB�'�b�'���'�2�'m�4��lX��̴,��(�K�7�"�'��'���'���'�R�'���-��� �ϕ)��t������'?��'���'�B�'���'�RMY����)�.P��<i��>=�b�'`��'>��'���'F�'��J E+*0�d#Ӯm������E�B�'+b�'�R�'1�'{"�'����4NyÄ�@5�d���X�)�'��'O��'tb�'�'#�g�43l��&�"b�2���VP��'v��'xr�')��' r�'Z"��&xܥ�̃�kV|u�M�Xr�'��'��'��'�T6��O���XT����,X�b�jq�#�öy��q�'@�Y�b>���&�G,��t�N��K����a�*A2z���Oz-oD��|��?Ac@T/T,�«7?G��s���?���~^��ܴ��$v>�������/O������R7F��`��� D b����fy�퓜er8�ʖ(H5΀Q�m��/g��ܴF�&M�<�����h��Κ� �\ܳW��+2g�Y{���r�,���O �	u}���$��b��f1O0�;wF�/����$�%Z�����<Ox扽�?�U-/��|��)���8���A3�E��F�sC����d*��֦͚�l"�!n'&��7��~���"�%f��?Y5R����۟�͓��D�6K�PXQG��A����;���xI��v�c>yA��'�����e}rӒ�	��n\�r#�)G�l-�'����"~�*�f��$���p��iu���Bg����4��x�'h�7�-�i>�!����������5j�q�����|�I�h��en�Z~25���ӀRg�9�-��e�'� UP�y�'�8�a�eB�(� �K��\I�n�r�'�9�gF�o]�\Z��D�h����L@�Upz(y�d�<bti�_9k�,t9�%��}x���A�|��E�GOG�I
��B�#�/JJv� ���}�Y�b��1~JZ(�g�(Uy8���&brM�f&�9f��a����i�H���?bYf��U�ĉ�R�#$�8R�N Ǣ�b��p��ʧ�0>�FF.rx!!�ω�N��}Za��v�<i���".��b�K�*z&��tl�p�R�c��,��`���A�Б���#3
�aZ�N� Rv<��o� iz��ӻLM��s�E�Rx$)��mj�#1����$��N�6�:b�ح`"Გ	�Q��A�톢5����	��Z�R���麰k���{	lXS㫅p���Cg��-l8ېn��|L�����2D���q�� 䜝��������C�	"wTLڇG��\i�}�烏7Z�B�	2U�-#T�
�(�1#�'&T�B䉷Q>�0���óU|��{�(��pE�B�	�G�����1l� �Kܔ!#�C�I�x�h�E.���A`$hբ�`C��2}��)�+P-O�P��1O,n�dC䉻SXj����'�qb�ΫN��B䉣'-:��b
���l�-֦B�ɲN;��$(C،�FN8}�B� NI����"��iO��DB�	>O�ꉙ&�_�=d�H�B�nv.B䉼�L5� Oއ&�ݘS�U7m�C���hE�s��4��4[pH	�C�	"` t�JG%[=
��(�&�-<C䉎6�b����H��s6͕5H� C�I!]�2����Q.�Sb�֓2RB�	��l��ȗ/4�	�֚��C�B5d}�(�7]3h	;���&D�C��	a�\ڱm½[r ֈ�Y)�B�	�Yˊ��A�u	˷�F�A`�B�ɚ[��U�N��c=Q��ȅ�C�	,��l؅�ɣR�4� @E���B�ɾ^Qf��S��&|�85�!� f�B�)� �0c4�Д�f���iL'	��y��"O�B��G� &��Jo�����"O��SV��nN�"��o=z5��"O�e+��՛ ���"C�ҝ 7R=�
�'�j9Эځ�0�w��YBpi�'���c�����$$5	0�Q�'��c��p��2IF�6����'N�t� �
#g��9���	2���
��m��u�4�ТU;�a��G�{�h�rg�S��d���!��e�|�*b'��|7�>�VrqZ|RB���b��(�O�rXaӮ�;m�F�i��%c �	�'p���1?MX�$E�Uz�u�'-����P�e�ReZ�OI7 �"r�C���,��Mָ~�|Њ���n�<Q�eD�s�B@a�DĖq�*�h��M	u�F;�'f�Dm�R��ܕ��O��H�0t�b��W��_��� @�'�J"A� =��iC��W�jX'LԀ9���h�+[�v�*sѡ���0>��FE�5��\�E�ߡk�tp���I_�'��Slz`�s�� ]�r�{�?���8��W�i:�s4؁yq"O��8uGY�V�c`E�}��ƾi'�)�˚� ��铤�Б=Q��q�t��5�!�$����4LV 6������ͩ�y�&2��M�d��Y�25��O�!��`#��lӘmq2F�F��h7\?M��:p0Ġ�����5�Ã�a~��Q+�Ԁ�Ղ�.5t�����+�����AZ�Y���PG�{����IE��EC�+U7��87�D�*#>	��Ù(�|�(�NͱYgF�r�P?q��/X�؝���4JzXh�&&D����"w%�(�&D���ti$Ji�,pS��/�4�B��Y�"��	���O�e6���(����3g$G$;N!�d��� �( *�sNx��ϲ>�&�����e:g��B/0�[ҏ,Fx�f�5"iT��e� \ۄH��B?�0?�T���ws��0��.���D��,}����ɬLs<��%H
�Ta}"��5>z���ɔTt�2C.�)ֈOD����W/1B<����=��d�Oܖ�H�a��~1Ն߇����'�rD+	&K
j9�s�^
u1�xڜ'4�a�����~G�RK��7�?1�#�Q	@��l��O�<���)0D�$�V���rP�@�bX��3"$�<�e̫!�2�	3Ƙ��0<�&���v�lK ��\��q� �pX���	% YD�Ҧ�ũ#N��84*�	Y��
���-_^��#��#��\~��u�6���)$�LDz�nR�Q��X��)�P��kpX4 8z�b�A�/!!�D�6��h���4#Z�#Ʈݯ	���M>v�9�=E�ܴWz��	�0sp�x����4��I�ȓ	�TI#g��\o`9�������'���x�'6��Q���Fς*6�B�q�춄��6OT��u�W�8��dQc�.=���"Or����/D�4!�΃&N)#��	�-���ق��*�:]����-m�r�k���=�B�I�jm.h��˺? ���M��6��%M3�a[���s�
cd�"�:EŻgD:���"O���@8HQ�)�LI�Y��_���D�
��e��ɝG��|ᒆ\�d]| �� #�$���� c $�{�|�ܕ�#��� �$��Q����B�	�V��a�� ^�D��pQg�R�V��'	���N�L`�AF���6�(� 1\q�� �j�Ӣ"O�ib��]F}�pTb�2��]�0�'o��R��J �??�Ϙ'��i���u�,�1�Ewd�0H�'4�k�GW�v��hP :nZ.|�rDT	%�t�4\�]���''�I���3s�jq�#� 3b��	�-E���R����uj�$I�V�b-L�!�4���ڒ\C�L+�'��0Up\ɲa�ffVQ"�O๐a�Ty�f �lo��D��c�0q� ܀��� ��i
���+�ymE:g{@��K�C0�u�vBC�����=�r����S���~�<Q��-0��;���"��L��) ^<Q�ˍF �0���#1��Qc���V²�oZyy��
�\��N���DQ=	ANa��\m �ej0.�axrS�/v�nԑ� Hp�L���d#'��U��B �i����	#�O�p�GQ�z̪G_{J$d����Q'����3|
�E¬O�+�L�?m�tM�^�u��fȨA��V�*D��$��M+PE��8���!Jh��۰
E�j����d��?�Q������Q:`�ᝡ[W��yf��[U�R����J���&7��ř�hq閼i���I{���:7�
n]�4��'q�n#<i!�2OW��S`'N�}��$�s�'&�x��e�"�M���r81i%�'/vQ�s�ʵx0 ��j�D�\t��j�}�]9�p������9Hq�AOAa�>�D��/R@�!nZ1TV����������<ͧpE����0����� �(\!��$�\�3�CD�@)9@�3'��@F�3�D��X�p�s8O��e���{���y7I-R���Q%BC[�����!���?a6g�$�58 �X�ZH�!�ɢ^v��fM�C���Y��c�V��S�H��#<�3���MH��� ;{��!R��D�'Ul@�$w��y���/�I@�~S��*viعzT��y�CKc&TE�3m�̦9S�Zt� I�cز\Y�����X8<&����ȧ>��L�-,D�dD����~��|��iA6;�J��r������P��K�<��b%S
� c�^������Q@5=O�t��IH~����y��W�p��:���,Nf�Y"�G����?���ˏ~a4�`�b:�����gSI��lB@G�)�~��'��84� "<�Q&��S*H��Y$�X�C�$�Z�'�t�PE*�56H"0
�"������h;l-�d�P�v�b2m�.]�	�m.��Dǃ��y��'S�s��а`�*m��I��B��%�Th��1��O��PĀ(�?�:`c��
�@�!�޴F7���#;0;��Ն
���Lip��<�����t���g��CEm՞b~\�jc�ߥD�B�h!�EB؟�J��ʊ}H
�[�σe�Q��8{I�����5��=Z�!�O��
Sj� 
���/����I��M��и<��"T��~ң�B;7��	�/ �Zy@	��M�<y #˾W����ə���;���q�;v��9p��쨟�hE�_�s�Y��S j����"OT8�
Q�q�<��Q�_K�m��C��������h��$��j��mK�ΆX�$a�� ��;�!�$�8R�;Y#�80f�¶)�"m ��`��1�'�VXڰX�5aJ\{$ W��Zۓ+�"�"1+�$� <�R��5�jl���VJ:!�$���x|�"�fX��*��ұO�H�-��|
��E��'��R��!�oػuV�t��j�ykP-y�0�F!�I��jX�41�������h��$^�Ԛ��f�Q�P���j��E�!�D  y�腡(U�� z`j�:4��	� )ҡ�
�>?B�	g`N;hGr� ��pӦ9�1M#t6O���F�
[3��c���FP�I�T"O6L+�KX�w��ع��6�H�J��I.��ɉ�鍮1��1{�cϐCP|� �*ӈK]!�B/AyˇNɼ� ����g��(X9Pb�"~n�2?�R��RF��py�	���72��C�ɻc*�K�h�R�L�"t,�^���{0�1a.-|O�Ԣqb�;:ԑ׆?Sۈx�7�'&��c���M��O�>HL
@i\�����vn�<�ä�4�&��"oI�qLnpJ���C�'o�bTD��H��� �H;��R�*�	eb��;U"O�H�fb�)v��\b	'J��p�i^��2�"�u�S��M�b��@^�,����T�L�h��x�<��`^��p��b�Z�Y��l�s}��W%k���ė�OI8<S��+@@�3wo�>h�a}b��v扞)b��
M�S�\<2��U�B�	�.�Bp�Z=_�p˧ �%+�#=YeU'�?��v�]5[u��`%�<��b�8D���:7����0���.9���w�@[��M�S��M{����&f�LȐ�Ӛ�4����n�<3�����%p�F�%CȂ�xƯ�k}�'��V����M�P6|}����}U���c,�dK�}b$�=�~��Y�d��G�Ҧ}��@2�y
� vq��rM*L�����Z��`�"O1���2T��(r�Z4f��Y��"O$p���E�6t�P�B-�l�#q"O��aW����]Ѥ�]2ZtF�aV"O.�`æ�(x�:h�,�fX9Ѥ"OPI�7
�!e�|���NHp���"O䝛ǭ�mT�;h�4[�8e��"O�,��јs��|Y�ś>ʸH`"O�Y�q��,[,�HG���tv"O�a����dal���D������"O��SH�;�~i@�f����'���R�XVh���gP�D��L��'Px��a�c0���g�/l�ER�'�>�J����tٙ�!�$���
�'G�=5/�9�eK�7
0k�']�=kd&3`�QEA�&e���'��:'D[-v���H.
t���'b`X�r�,<FX�ABړU8Z!��'����Q�N��I��h��_!pt�
�'XЈ�&�/%Ҋ�QHɯW( ���'�����e��I`c�JH�u��'��4���� u�Θ�d+K:	��'30�7'�).���^�1Q�}h�'�<��5�ӞB�"�x��-xR6"Oᓑș�r�kFڡ�i�"O��܍nix̉1�|`#a"O6-S&*ə0x`����?`�PI%"O qx���
e�	1��;W�EZ "Oڅ�׬�7W�����6U�%c�"O� R�7�@�B�n��،"O���n�6�4��-ۉ>�b�	r"O���I_�4��]�m� =�ڰٗ"O 
$!��*hj��H�S3V��"O�=�X���Z$Y���3"O�A��E�/��:((n�Zq"OT�@w���w�-p�X��bM>0X!��@6�P���-��՘c��+bI!��^�C�F���
�]��в	�!�d�3bК�S`bX43�$|��͊!�Ď= p��T���g��P����!��I����+pj�w�`EaLZ0g(!�GP����"R<fiT�K�(��&!����6��$Ό/��4a�>)�!�B/(O��k`�������!�_��P�h��Pd�t ��Ь/!�d��	e�M��-^�>S�8zvj�	�!��O3Ծ�����8FԀ��K�-	!�!��\��	֎>���H>M�!�Z({T��:��ˤ(� 2�A�!�dQ�o.���ݞ<=T���d���!��/i-�uP�˖)�Z(J��W�!��Bs^v��%/	+#��r��k�!���$툴�De�2#&��5j��r�!��& �}�3딓F����&�,�!��ڞRb�쑖�H(t�`����`!��+_�@��[�Fgd��CU�6�!���0�2`��a�8y閉1c !�$X�*��H�s�_�Pr�U�� �r!�d^]LPR%��x�b#�.��?�!�ė%)N:���%H:�|�U@� 5!򄃮o:Μ�@`�2G��~�\�'����O=&��&�I����'}�	��aU8C�@�xF�{��%��"O&U�����G�l*P,�#* �A"O� DMh�F�Z`i(���J�I�@"O�p%ʌl��M��F[��1"O$��-�*$�Z�h�)c?hux"Oh0*�@_�<�f��塎�6Re�#"O\��b�-{���Ч��G��Ћ5"O,�S��T<4\�y! ǻK�D��&"Oڅ� �T|@�/�#Y��l�u"O�KcV�ml�`�:/��4Z�"O��q�� �ƕ0��vyޔ�"O@#S�Ϩ�@)��>c=���"O�p(F��u>�IA���;|4�"O�xе"��+�0��ُ�Э��"O�}�5��J�NHxg▣a즜��"O"4�E�*Q�F��� ���	�"O�Aw�V�f�6�P�+�����"O��@&��9���@��b�(bF"O� ���Y�n�  ۨ=VJQ�!"O�y1�gT�cT�� �v>,��"O@9zƣ�aTP�����Œ7"O��V�S�x�z�BE��4��p�"OJ����b�N�'+�0�┚�"Oʄ�����b�t�gi
�z�nQS&"O��M���R��W���|�,P�"O�m�gn?|���B䇷l��p"O ����7��fC�0i�x(��"O�$2��֤kNܱ�� Kh�qkA"OZ��.�9혭�� N�]:c�"O29Q'�]�Xy�E�`5�"Oxd������$D����<}p\8"OؚU�-�{W䒎6|v���"O|@rw��!6��3CS�o����g"O�)���0\�ɨ�O�]ap"O,�z��ܦU��,��ȋ{�n���"OB�x��E3 Q��U����`"O��R�G.i������+0�5��"O�����/%#�x@���),<~���"O���t'�>!\ ��9a�ۗ"Or��V�E�����6/��"O�A���T"h�q#�6�%��"O�����E1#!^�7�fp"�"O��;���iQ�M`a�ղP@q"Oza�`�W��D˂�F�S�8�6"O�5#�6��4Hb'�=?D��"O����J�Z��Ʒp>�l@"OȅB4�ҍL"�I� ֝8�T�"Ol�%F�L�����nS� p� u"O��ҠL2v�<xJ0K��$<̳@"O�!��K-J/��b�)N P�r"O����d@���IxǇ�>' #"O�H"4iԚ.�0�2�fC�r��`�Q"OJ	c�ˏ����p�[-lԎ�h�"O*�S1�ŧL�~ �bؗ3��=C�"Ox1��O��_{.P���ڴt��ѻ"O,8�`�XP�C'�
�g���"OR͋�B�>x��!��4�f���'-���ԮS+ �p��4ɆQo�I�' �5p�G&+�4�d- }�tB�'� �jc�݁W,}�����x�lu3�'�@�&�#a�Լ9$f�wF2qZ�'�t���ہ ��Pc�ov�`���'���C̋*�2Xin�oPT\��'�xy�C,]6.�R)�qf�3?����'z�x:RL�7'�i�g(Ķ&'����'C.�r�B�tyw`�i��a��� BE��N��m^74˖��*O�5ӥ�ˇ[K���`خd\<̩�'�zႄ��<�h'�T'[e�mb�'��-zC�E�k�d8�VĘ�_Rk
�'o��R�^1G�6\�&��R��'M�@+uE��D���&�"p!
�' �)�M�7Z�d�X�h FŶ��'������=m�R5	�/r&���	�'�8��Ӯg�p�P�_�kJ2��
�' �=��A��va���éQ��dP�'�B��ٝM*�$2`B��(��'_"��d�ֿ#p�t�'�^��Yi�'pXqї��$N�`����V�@�'<���,�"\�rؓ ڐ-!�=��'4\<��g
�DɈ��)��OoD�P�'�$����\�K��M��:����'\\����O��=��$T��n��'ݒ�y����R���5@���!�'#N�j�n�O��@��,�rd��'�t�c�S�QD�A��L�V��P�'���@EO��Q��U`�K�x��
�'A��
B���B垭V] ��'ӆPZ2�}E�I�L��\="	�'�x���׬�by�en6����'���"���(I���'�Hi�	�'K�-�e��ra��
 @j��0	�'O����N�T��C��7@ eA�'.���tG�3.?y�딛�uS�'�*�A�A#y�)'��:~�"}��' �T��ܶ	`���^�*1.m�	�'S<�Q��'@n(���l@�5B�'�����L�#ˎͺ@L c՘<`�'���S�ʪ�,�{`	Y^in�8�'Nb���䛔L�@���n�2[�2�'I���+}C>�z0f�)kR�d��'�­,�=��i�" PX�<�'�� 	�M-}��	��^.5ʶu��'{��AS��,�LY Ύ7��t�'H�i«��z�V 1�x���'���˕ޗ6(��s�V&?fF�9�'���#Gʘ:�L�Ci2�\�H�'�Ґ�dh4zp��R�"U��I��'��Re��M�p!u��< :
�'�5S�E=V���C�	 �l]Y	�'��5�D�5_,p��ʓ�4)	�'i���� �G�8�X"+�:]Ĉ��'� TY��+f�v\�Q�^�N�D��'�YzVY_I��*���
}��u��'��C4-A�B�h�� �y�����'���۱M��.���RIP6�a1�'�d�Z#��?SH� ��U3�4dY�'ӊ���W`�<��1�N_����'%���@�P�H��8�ʍjR���'�hyxSo�}8���ޔo�8��'I�9C��V�M�4q#Ю2���'�l������GhJ��l�&�1��'5,���@�0�`�afFޕ[�� �'&�$�S��T�☀��S:)O`h!�'y�##�t���@F���W� �'1��b�-��%0A1㤆5W�̹��'�����o.%������6K�<��'���A������K�a�>C�����'|�Q��վI8�ae-Q�
�'��P*��L�B�ȯ&Xf���ô�y
� ��
�J�6O<<�A�30�qD"O�EK@KЊtn��Y6-H�X��\� "On���R�XDt*2L��(R�	0�"O�]�b�G�rEN	׫�>8���"O�x�B@�1o��P#�ѫr�"03�"On�'�#rpڅ�f�˿k���c4"O���F���:4��ɐ2�dq/�!���(x֌,p2
	obuxq�2X�!�ē.U��H�B��m(�ቄoS�B!��P9K�@��V�Q^z�Y$!�� �!��%g�uJ��K�`��,a2��!�DP3J� �*N
{�X�BnP1?�!�$�\�i��]�}�8�ycك`�!���Z9��)�<(�V�#F�[�!��ijzY�!�� �̈藠͌p!�$Ɲa� (���цu�`����מA'!�C4�y�2�߲!��A�r��-w!��S!}��$6 H��B,Rƍ�_!�ڬx��A�r@P�%w��y���F�!��A2`Y�C\WR<(ᩉ�_�!�L��yv�ěHr��v�!�����&�ϞkB4��2)>Q�!�d�"�����yR���.����'��jM� ��]9aC���@�c�'8�H��'Ҽn�"�sS��*}8xz�'�D�rSȝw��I��@�HiJ���'�Cgbճ&V�AJ�d�j��i!�'��i���7~��Ќ�?d��б�'#����>�	�$�ܴZ7YR�'�jL����Hj��g����'J�b"+K�S��!;�*ѿb�^��'*vaB�?Q�tbwѨ�F��
�'jᘰ�ƥhwh���-ƢW�t��'ƪ	��ՇOph�+g��$TL�1��';��Qo@�+�)����"�p��']�x�"kQ�t�2Mz����-�3�'�*\+���'��ؚ�d	r�40�'{28��"[,�[f)F ~�A
�'�4�aᇅ+�����h����'�l�q��V�P��SbM�(!��'�:@3Ƈ�C+ ��H��X�1��'�Y`�.\rh���.U�����'��T��LA
K:�r�M�d���'�"}� m��BP] $�I;pmY�'�$��nx����K�O���
�'��Y�gB�C�l8�c�:��
�'��C���rM����0�	�'W�ܨ0M'"|mH��� K���'\>e�W�O>:�X0� !q��[�'hЙsU ��@�*]�".U h�d���'�sw�va�염}c�a{�NP9�y��UL<�3�O
o�52G���y����?BhP�׬�gc���3�y�"=�(��Ja$��!DD1�yb;�Ht��0%p�\�A��6�y�ϋX���+u��R�L5Z�H��y҄�N���$��*K�-���Y�y"��<�NL��!:�)�v/W��yr�	Ln��̈́(:1Z&+�yb��$x� �@�6�����ͭ�y� �?|%(ŌI��M�#LL��y�Ç'V9��� >5��e���8�yb�I�nW�3�倒1�5�����yROO1;}��8BΝ�#��ٴjϛ�y
� ��1c�*E�L����(I'��$"ON�Qp'�` ���m�}08IJ�"O�*�H��/� 詆Ʉ.�%	�"Ol�8�A�<M�6��̊�>Jr�rA"OxA�N�"5>`U��k�e�lp�"O
P���:>�6eY�I@'U�8kd"O����y������` �u�"O�h�Ϣf��p�Dr�2-��"O�]ɡ���p3d��k�b �e"O�I�Q��1��Iwb0v���"O�y�J�!R� �A!CW�zeX��"O�p
��Їc�c���tN�(�4"O�58�E����ī
m/eK�"Oچ�ĕ!��E��#B&"��h"O>e��Q�Z�zQ�7���"O�)@'�w�81C���+���"O2�hgFX#���w��"�P���"O�9�T��`�N ���:;�
4iP"Obe�		dAr�@#'�U+p�#"ONX�(͚-�`	�L*-~�l!3"Ov�z§�R�vx�+L�v\*Xt"O�Q���r4�K�L �p���T"O���S������K��W��]�`"O��p�B�,<�b�ː���`��"O���C�O�$�k�ʖ�0%�ݪT"O����ڠxL�@�ƒ$H�=;!"O���l��%�Τ�Q�}��1��"On��玆*�d�Y%i��V�����"O�P�U
�VL(qHZ?>����a"O6a��B�c��܈�f��j,��"O� K��Y���j��8��Q""OF`��!�5:�� �]�'�B� "Om	��D4 8J�e � BiH��g"OzȔ��
�hC�O�d�`"O�U{��WJ�&=��-KZP��˷"OEhE٤?����g�ڃ"�� 3"O�u�r�N� %�eA$q�]��"O8g�ڨ
b�q���zb�9{!"O2�km0��Y��Z�ư��"OTkBl�"5et9+S퐃=�h��"O�ٻs� ���i�̏8����"O6�2��ڸ%}��+^��T�Y�<A�.J����&�$m�Ұ���PS�<����K�z2�Fzn��&�X�<A0�V
����N�����W�Y_�<�cu�8`�힀$��-�	�t�<0NT�sW��`�#ٗ7�(�t�Fp�<qv�^4I������^T�񣤉V�<ф�jCr�X3G�<'�xM)WS�<�u-݀,`l<s��6S��0#ʙO�<����̣r��>\*)�rD�<m� ���UA�?R&���aYK�<)����X:�L�AT��扙�OL�<�1'Ā��=�Q! 9%��m�A�@�<AS��	c$�x�/	 C�$dQc��V�<Y�A*6���@5�J�"����l�G�<�7 B23�|ȁ!��~'�]{��G�<!�Bi,�1	*��S�h�<�@I$t/H��S�·*�ԩ�nC|�<�.�54����E3q�����z�<�5g��|y�n�33zT�,Y_�<��e���$��� �?*\�7/[Z�<yQĞGJ��@���,<P4�"aC�V�<��I�+	g;�*P�x����7��T�<� 
�y�ĝ;t=r��0�X���q*T"OM÷C�J�*}�I��6r�}�u"O�M�WO�5�j@b�<Yad�"Oh���@D�BE+ШÔu:`��&"O(�Z)��C"cS�*"��&�y�<���E#���R�����)v�w�<AW�ڃ7V�j�����Yv�<�1�dq�IF&�~�Tц��G�<��@/06ݺ�d�m`�3�BY@�<�Fb�s @��D���
� �y�<����49΄�G>,�m�t�<��g�I�ƭs�(�t3����@�j�<�^� H��kgC�fe�4����d�<97���Uʨ�	1�BpBz0YQK�k�<�r��r�|i���=�0�ca��S�<�#�R����	;�Lġ�Ǎh�<��D6���ҔL[*��t�2�O�<�b"�6+xA2Q/'y<���a�<�A茾{�u:�K�3w�̀�h�<��i��|���(��D��(XC�A|�<i�e��:k�2�+ ���ţ�f�@�<A&�"l^�Q	vo��h�@�c��T�<�sϘ�a3�	�K��ui�����RI�<��eS�B�� �b�20<������<iR@�3d�p�p��B�)�|��Y~�<As!X��=���U:6��dK��TT�<ipf�5qJ�0êH3;frh�w/E�<����&���,M�iW&�hcJ�g�<����):�f}�$*�{�*æ�`�<)E��-~��3��A��.Ѫ�`^�<� �4���i$"F�D�W.\�<��Fsюt����#z΄�dD�Z�<��F%��P��� ��X�<�thN�jg�Ѐè�r��%3�!JZ�<����$%�<<�q�XI���C�z�<�Ҙd�������#Y�)�u�y�<AS�J�=�T� $�I�.y<��F�s�<��AWr� ��?�N���i�<�lX�;�0U)�gN.]��M�<	���l�.LS���u��b@-�J�<G�ӂi�K,o�5W�O5��C�	�)�J� :��\�5�Z`�C�I�Djh4��[�uT���g�RC�UKj��o_,YT @��(|V�B�Ɉ3j�9���B!	��ps��PB�ɨVC�ԉ�H%��p�M��$B�	w�>�Ӡ�Ƙ]hv��ă�7��B�ɑ1���e��#�F���	�+g|�B䉁&_��;3f�0y�.�HQ*�;®B�	�o���9��N������!D'!�DɲUD����)��<��`�!�D�dr|r�� �����*��!�B�uѦb�UxŲ����J�!�$S ���G�L�r��V	�!�䕉�¶��/Li\�q΂K�!�+fw��"��	T��%�N�!��I&!�����!�!�d��R�!��Z'd��ЇQ�jxdW��9�!�D�'�x C�c��[�ف�O�2?�!򤁽�䔃�6'S=8 ��!L!�D�\�khG?�샴��!��٭<dX�ڷi_m\JD��KK;:�!��|����oQ�k��-��I��!��	$U�J4���ùj3j�[�WG�!�� T�Qe�b�8�1��V�Pw"O���B�)�Шp`!ɓ����"O9�"n��7� �Bb�	l��U��"O����ֈ0ʙ*���2�X�0�"O�m˖���Ux�4�_=�[�"O ����*F��YpdN�h&~�r�"O�-�U@"|�)���� �xy�'"Ov� `M�v�`�%s�*	�"O�}���|3"-�@�8��x��"O2�% P�K5+��� `�� ��'�ĝ�E`�;(^�x�'쓀��L�'p����N�byĤGj��R\��0�'�0U{�F62���#�͈E�d�1�'}����U3m%h�p��7�p��ʓe="(iGÄ�nQ��{ �4-Ѕ�3j�R���1Ϊd�dʞ�( ��^���
�ǘ�z���`��#ֺQ�ȓ`;�����Uj��0�b���p���Z�B4��3�"�&U31P\؅����lܣ�Ɓ)p,�	9�H�ȓ^2PD���$/����������o��m��ԵSt�M�@�*��@�ȓ�*y�6�^Q6h0w#� Q��A�8�3,	]�6P�+�+��A��:�Fy1� �7��s�J�2 ��r�4�FFɆq9���@�} �ȓt��M�T"͞
T s�,Y��܄ȓ}SR\2�T��p=��׀D�0��ȓ)����V�,<2�I�Agҹ@��M���L,�G�,�R8���32+����"�K�����k�P&ml����'U����ITHz��)@70ͅȓrp��."iލ���ؠ��ȓap����]� ߒy%� ��5��Z
�&�@q�E����s��ȓrP��g��9,���p70*:.]�ȓ@{\	K��0[����'��2~d�Ɇ�B?�Aۦ�Ǣi��8�B�;xp�ȓ�
�:FN.��=�ы$r���ȓ[w�5"p��"�B	��m�Ux�x��pi�hR��^>��R�]���1�ȓW��rP��*���#6��54�¬�ȓ ����A٢F� �����H�^D�ȓYl�d��*�N��������ʓik����l�Q�|�&�6zQ�C��m�2!#�gR6L ��;�#��^*�B�	1{�,���VI�@��c�|�nB�ɝ
]�$(1�Z�,KL]�c��dB�	�Nw>��yr�kFAߛ}�B�6Hj&�2E�y��9S͛!rC�B��10��*�L�!�����Γu}VB�	(F����%Ü�~�ы���%	�B� �l5Cc�+@�2�#��*!�C䉃 ��tʍ�0�Jd����>b�C�I�>��M;�kR�:���*EoN*@�~C�	�#�b��F��1L%~S�'�*EuzC�I�UB�)�g��h�8c1j��A�>C�IhbE1���&O|-�����*C�I�Oz� W
�<eB�t��ԣ
T�B�I(aJT�;��OW�@�`���^sC䉼crJ0(2b���f/ΉMբB�<WR*�!�NP�� e�ԫH�q6�B䉅h��)D�޼Z6��eE�	�B�%{�MI����Tj��V�-IhB�)� �)�ԩ ���@��#=�bR�"O0tc�F�d�P��"E�0J���R"O����nU?Wwj�� �]�< �C"O̬��D.$��#"�qNH�G"O�H��aٲd�X��Q�Q�^g �Y"O�%�ĦԬb���*`�K�I5VQp#"ON03�o����,�6SI��"O�|B��;?~:�f@'f�@�"O��"X�*�
��`f\/S�a�0"O ��&����@�E\��"O�� �K?����OҰ� �v"O����c<.�p�L�y$�"ON��D�[�N��sьͨN�98�"OB̂$�Z\�5RW�׽,�0�"O�� �32���*�mKt�*��"O�#�M�5>��,A0%.zz!�$�
#�@HG�_�B�6+󂎲!�03������A��Bp��9L!�D�"6o��&!�<q@�����k !�d�3f�ܓ���#>@�I��
�t�!�$����IVjNb��x�d�E� �!��Z)!Q�ؗGp ���M'P!��t�&A���P�ǹV��R !򤉑�b�*� �� Ul�)�#%W!�$ō�~pل�ە7bʬ��j�?uG!�$��z�×�/M`(`w�2t!�Dх�lY�*G�v;(�s0l�+z!�&d��s���-s.����! ��!�$�02�����)�9	v��bq!�dU�@4E˖�ӱ,��E���_!�d\:	1RA*�.�&�*�K�
.W!�U�DC^8ǃݡQʄ��!��*XH!�B�`�(��큿b�RӤ��"N�!�ĈGse�J��m���X�B =l!�dd�4(ǳq�
�d�Rl!�$�:*g��櫐7Az2� ��	�S!�dY�ZϒŠ�ֶtj�P �
O�!�d��X7����b	X5��v�!�ç�ȑ񎒴���K6!�!��?#�D�r�iP/��z� �:3�!��#+6���b��&$�MKՄ�)t!��ɔ|�Ȕ��A`$@��*bu!��)[M<�1N �t%X���"5�!���	���igܕp�A${�!�
�EV��&�_�O�ܩB�f�(k!����*��@$�*0Y��G+.a!�E�u�\��-�z������ )h!�dO~�Fu�!V� |�2�bW�{�!򤞦]9���$�'`V �@�^�p!�dǣ����r&13��)�E �d:!�=����E�`��%	 E^G!�$�$CV*�)H���@ �k!�D�Ig�x��a�%`�e��K� �!��uCR,)`�\9S��8�)�!��2���ա]Eּ#V��9K�!�ݹ\=���P�ցX2~*SA�{�!�d� in�����5�����\�!�^9]�v�� �?0�	#d�[��!�R�<s��ɗ��:R�ȥBf�~�!�Đ�Bb�8�B�=��-A��-u�!��4xJ�����+}�*a�@��5(!�d�f �Gk�� h�g)��Wn!���A�����%F�>� �I!�d�	g��Y��Lr�ji�Ҩĵ<�!�� 2��u�UtU�����&>r���T"O�X!î?N�Ř&�iAt�d"O������aXưS�L��OP`@�"O)C�=�"}1�BK�C�� zE"OHU��W'"�k""��b|��[�"O�ĩ��_/$Yjp8g��bɨ5"OV�闆�*&ډg���?A �:"O�r��R<��e
�2;����"OL�
Ŭ�/<���S�	,9,q�E"Oa�T)f���I�RE J��7"OtQ ���ey<�2�'�4��"O��&Ćb��;2���y��"O�A�猉*,�� �kpع�"O*��'B�ۤ�P�O)ER@! 6"O! @Æ�;s�VJX(%"O�����*D�ݩd�;	���y�"O�$Ц��qJ��j&A Ԥ�i�"OfYHabзc�pHƊ���qL#D���Y::=葎Q�d/��2�3D�l�� jv���E��b�H4.2D�l�R�͖T��Iz
[q&9R4�.D�H�Q�J:U�D�����}$��K�+D� !&`T��<�p�^)Wxh4f7D��R$[% è=�tf�4 �,����3D���5+Ū`��S��Ӌ|���Ee3D�X�A�|������p��t�$D����$(0��Wi�6�����#D��$Y�>E�y`�l�;w�~Q	�j+D�����R9Na�Yxt��*wG\ib6G6D����M��+z�{�.�u�.-s�4D����B�1ؾLm�9���1���c�<�v�X K��9 �1>Cր9�c�<��̔}��ܘaD��<�|�T[�<�eD�6	�$��6��U��X��s�<�V�]W��D	�.y8���c�<!���9&�)��&AI ��5�Jv�<�2�ţ:¤3E!��Bښ�8��t�<a"E�Z!���bKT�~�tC�	0V ���5��b�"U�A�bl�C��?~h �j&�Vl�wM�#7�C�ɛvތ�i2�Q$ � dC ���C��:}�Hr��3n��<2��߮R``C��/+�R�s��1�Fes�o�"=�hB䉓6��]�3L�d���A@Aq4B�	!C��8�Sm���0C��B�	QӜ�兛�slT䳔��R��C�3D�ƨ��#V8u�4���E��C�	t.X�!�o<Q� ����C�5g~��h'ES2�Z�V��B�	�(K>`%4D&-yV�'�B�	�Z,�t;CJ�7H1��[B �/L�B䉐H�����^���a��`��B��;%�@I�O�M�B�)� ���B�Ik"jh{��${Ʊ��@�%�BB�}�l��ծ�.�n��F�QB�ɱrȐj/�,����P��rAA?D�`(uKS�dzډ��IE�`�o9D�p�V��aPR���h�v_x��8D���C�7�^�I�N'P�p$r!g0D��:׍�\���0���h�d�a�"D�����,|
TY�R�	� ]d����?D��1��6�J��%��!�F8�h3D�Ј�N� �����n*�p�,D�lK�/;�l�����!��a9�+D�� ���X�$�K��/@A@���"O���ǘ".a�L;V]�],�!ʃ"O~Ec�lS�4��1�	,��"O����0�� wB�Z� ��"O�D����I.�t�0���|}��"O��:�&�93�r�!���c��l"OT�ꖡKX������J2"O�ĸ��ɱl����Kݍ@B,��"O`ݛ��Ɲ_�`ۀ(�_CPY""O�8�L�?w>���&''  �"O��S��]=3���F����M��"OnA�����P_ )��Fħ>�lR�"O
\���N�ei�Y7��WpZ	�"O���AJfa�e(���Y[�q�A"Op��K=hTB%P`�!I��i�"OXy��G�z`�ٿT�^4��"O�V��J�!f��AM"	�n�<�d$ɰš�&�a0����Ho�<Q�E]4� ����G�u���j�<�P �>2O&( �[�qz<zg�Yc�<�c�
"}*�){w	
7'Ҩ+��`�<���W�nj�� A� h9fQ����g�<�a������@��v�C&��j�<1��	�^y2��K���2Efn�<Q�JB����!	�5� ��w�Si�<����1�J�e� O�
�;0o|�<�1���9e��0��ס��a�x�<9q�޻<8jty��֩R���'��v�<i��űy-l�zNC'd���x��I�<�I|�t �n�TX:��C�<y���t#	�`G�75��8S��G�<1��O�IМ$�'��'�����IB�<qUD�qD�q3�b�9
cvT���H�<��á0�h��U*Y80�\}�2C�G�<Yw��!u�5:�!K�4��˰(�o�<�G,�f��DRSN6-u�1#Q�<�­��t�69����1lGu�<�R,�%}�X�'���@;󏅾�y"k��r.��O�Q��H�qa���y�E�5X����ؔ:����I��y"�R� ���j֘b��y�#�yr�� LE��"V�ԽR,��cI5�y��%'7��`k�w
h��Ua9�yb�͜V��Չ[ ��I�2��y�޲l�8�`����dU!��̽�y�N�4��W(�nwl���C�(�yBJ@�R"���O��`.�c!L��y"��V�`h��A�ZA�@r�)�0�y��]�4��8��ɭR��Z�"/�yG��z�Q'��tt�8R�lC��y�n��E�`2� ����r,���y�AL�_����r�׉�8`(Q�
+�y����
u!�P�D��'�ޕ��^�>���a��C�`���'P��3���k������'��������=��&G�X��d�
�'����H�9�QX,�;��
�'
BQ�Vb�
Hh��	(&�PI
�'5L��s�/|�*�	Ӄ�$#�P�	�'9�y"q�L��~A�ʂm�Ђ	�'���2�] �ư ס��j6����'��A���)Z�� !�̘ь��'�a�Q���P�eѳn�Y�'�� pր��qL�I� I#��r��� ��v�=SnVxI��B�f_n]�T"O8�څ�2r�����cyf��"OR�f�4j6W���(h�U�O�<Y���4s�L�;���DE���YH�<$��G��H�cBйar=�C�<��S� [��A%�U[,��� g�<i���`aV ���  NN��z�<���0\Y�iP!Ȼs���G�x�<Y��1�|z5D�5"��#EGx�<9�'�Yh�ȫЫ��k��ɣa�y�<	�o��y�CA�_����L�q�<��eODhl��3	��B%8u!Bq�<��g]�S��0�	�<&0x{�G�<�u�\�u$�B��J�B�:=��^G�<��O>ܺ������	RƝ��!�A�<o@�k���f�UM�<�S�<Y�ኙ
�-�u�X�|�r�����Z�<�Td�/C��! d��/�d<�p�EW�<	��_�7��X�h <u$f�	U�U�<��L��`��t/F�df���7%�k�<!� ��,ಕ��%��D���A��r�<1�,�K��� bA�a�ębw�l�<��c�d�[���n�\@B0B�r�<��Պfl��	g�]�Y|��
f�<�&�D�0s����F��oJ�u�'�b�<9cH!dչ��ы7Δ�k��E�<�C�G��PHu�H�a��I�<�G
�3x/�q�	7 $��b�B�I�<�" �rE��:͝�/�!"�E�D�<1�h׼j]9D�?�� }�<���
� ���P"j�9���B�<�q�@r���+L�-�܉iF�Y�<)���X	��m�$���1�+ZR�<�PC�&`[���M#h@��Q�<	�l	�b]�D��Ls��RO�<��
C �89�G�:�hE�<�bK&[j�I�۲8����}�<�n+nxޕ���_/4B�l�|�<���Fn�S�)�,�R$�x�<�F2v�u#�X9h�\��fF�m�<1bN� �줒q/�<!@�A`��c�<9�(�
zl{��P9Z��T�I�<���מ`�\��F�A!N��uC�mO�<���!iٴ�p�A(���B���C�<!��"!��I7A� �:Q:���G�<�#"�<UԼꅎÐ�豔dC�<�C1,x�BU�6�thWe�{�<頃 �4XQm�=DR5��z�<� �W���"�ΥKi��!gD�P�<yJ�9=e�� &�Q�6$f��7!D�I@��,1���hR�B�t�j	) �>D�,pAa�t1��TK� �hU��=D�H��"h~�b�$G#-�8u;��=D����U�]�ap��0#�&�'�;D���V�����p���� ٫78D�����W<.g�)S�)\GR���&7D�`Z�	���fM�� ۲�u�	0D���#U]�"%�Q`�0���o.D���F�X(E�$���"�m��ka2D�(y�d�;��m;to[�e��@G%D�DC�ő�]l x��^��R )D���b��eR����˜R[�$
��$D�D!��'�rH��ȇ�&��PrԎ/D�"���NQ��K�d�*��"D�� ��D�ʕ	3Z�� ��k#�� "O|=�c��53��(C�]����#c"Oʁ"'���eS��൩�O����"OZ@�l %������]K�e@`"O�m��B����r���
&h�"O����ȕ�;����o��.���"O��$�j�~�AH[�[��dX�"OhÄ�.�*0Rq!I(Č)ӡ"O�|(A�V.LZPY��	.S�!�"O�D�� $�a8���!�9�"O�Q��N�5^r!4��� �0X@"O�5
ƪ5��8HX�$�N�b"O���ц�(UFI�GS�P����p"O�]���M�\� 4����2���"O搘rA�5%H�&�у���*t"OQ��BQ .!`��� Y�X��CG"OVh+ANp���ʓ1l�%��"Odܸ��&9c�!���ڀRH)p"O�i��� a7���`���M= ��v"O
����;*´�WN]�g74���"O ��L�;C���MA�X.�ش"OĘ���P?Ct0`�,? 6��"O|Q�B��9�<����*G ���"O�%��F�!�vը�D:@���"O����VID"H�j��L���!"Ov9	��[�w�~�w*�+��䊅"Ox���ճ[�j��B*ֵ$|�)C"O�2�EĈ������^f�pJ�"Ohe�Pk

H�f1����=\aN�t"O��-'8Br5��C�v�6�"O(d�wb^3Uj6y�V)����"O��k�(֟)P�"p��h	@W"O�-��EX�xn|�uoݹa�(�"O�X�v%�l�X:2�X�YZ�C"O�pt��/��M�	׏}v���S"O@��sɝ�	�@D�4��we�]�q"O�cD��t8�m�C'֋2^�Q�"ON,��@,ws.�@	�#fV�X��"OD9�@ ٓ/r|!�a�q8R�4"O
��K@
	�V��2��$"�y��"O�t9`鍻vg�A;���>��0"O4Q���4.D���܄L���"O�=ktژC��Р��)9@���"ON ������Bb��"EG0�
�"OġAa�
7$`pM*��E�@�q%"O6�H$��6Y���!HV��1+C"O�D�+f�C��!p}�|ce"O~�ca�؁[�>U��
�Uon$,�yRA��bXi@D\bL�$ʉ�y���$�X�Fd�[�>��2bZ��yb��,�gB�5V&��*"���yBi�����UdXe�%r�'߇�y�� �� ���I�ک� ,Ʈ�y���*}Ϝ�R�ȏT6��&�Q��y"k�D`��j�F��A�`˗�y"U����K��9N,:�	!�y��ڴnxF�j��6�����y���(r�d�2�A7���U��y���&�0<�j�4��]:Վ�'�yҌ;,`T�&H�&}�����ء�y��[�O��a�AR4XH̑�B��y��;p���	��ј[ޚH`Iҝ�yb�
]�VF�[���R d��y�/���\�A�Ou����R�y
� ��"$�NV�����u=M�u"O��ٰ@j��$�EJ�3\Jɩ�"O�x�$���/Pr@�wh�tOV� �"O�P��%/!�DY��C�fC�]�Q"O����.�%:�.	��΍k*�U�T"O �4��.{؍�̖~(���u"ON=���MY��D�6��`�Ш��"On��qk(`�������OEXAxd"Op8J�)|�(����;>�+�"O(5�0���hq�䙄U:��:�"OHA���)���hve[$h`x"O��HE��^�X�j�;q�����"O���n�y$iB�	ʬ�V�p�"O�ųÁ�Y ��
��^�1���!"O�(��ߦ%���sg�$4x��R�"O�)J�kG"	�P��A5Z�h��"O�Y���)��ɛ0��_Rl1�"OV�#���:���%E\BݼD��"O���%-ߓ�h��J;*���$"O2��#㜜fhe�C	�1B��)�"O.��2��z\D�UG�b'�Ȫ�"O`��3L�+O� pL^h7����"O��pd�޵)��U��K*@��0"OF����K#o�ZL�sŇ= Y.���"O�бp�a�b�A��D�.Sh�b"O�АT���`����/{q�P�"OF(IPm��:����BO-sL`��"O�xP�΂�d��f��U�) W"O�be)<��!:�$R�J�!9u"O�����?Ih�@�CZ?S@D�k2"OL�v��!r>�ц`ȁ�~�s�"Od!
�O::�#�/�(Ōi��"O&Q{3.[1���X��U	,�� �"O��$"�|"~i��צ$�r�h!"O H!��V� ����,z�2UC�"O�hׇ֠i���t�[lp�'"O��X��π[\�=�6@l	aahL*�y2�WH6:5��B1|�Q ��ybD3C/u�0��u���#m?�yR�Z�d��E���W�l������yB%D%4;���_/v���Ö�y�V������lH?O1<q(� (�y� �/ ݮ���䚬J� ���<�y��^� 	�D�v/>>l�X�#�J��yB� ]מ��\Es����*	�C䉺Zf�uRR�X%|�х-K!
�C�ɵ4N�PtM2<��XSA��D��B�ɲ7O|�JA�׮��f�k�B�I3*�T E͘M�0!���3N~B��&r�h]�!��zchx���gFB�	 3�� 9��*2��x!�A�W�
B�'D��m��o�uf��(C�.�0C�	�M����Q��Ee�R�K	{C�IhH|�����՘�F�m
�B�ɾAd��O�V�DY�X&�I��'	����Rwv-�$|�j��'k�<xS2;ıc��΅r��i+�'g<���L�4ܝ�!b �3Y#�'��R�T:�(B�N%/qV|R�'�Y*3�	�|V��P�P()����?9X�$��a�p�0H�~/�D��]��	�5 V$z��x���T�N�z���M�ؤbDBB�RX��Z���� D'D��t���0�p��a�RD�#	$D�� ���hT.#�(�H�I�h�Bp"O8	r�KԧN϶����%R����@"O�q�'�mu%��$Q�KG"O�И j��	����Bպ8ڜ��t"O�aP�!D/,�`MI���.���"O18�-N�x����D�O���"OB�I7���tД�0v+�3:Px'"Od|�Du�2��������"O\�5�]R�2l�@�_�ʨё"O��t���wp�޹N�>�� "O*Ecy#h�S�
\}�Е��"O���g�7�
�[@��m�.�0�"O��
�@����@AA�q��m�r"O��B���b���aϪ��$Ѳ"O��*��Q"7)H�C�ԝyp�y�"O(�����&wtؖ*|I2F"O�tR�+SYU�����!���4"O��iv�PT�>�I"g�#��)�"OT����Ne���r� P��Mh"O~tAf�'&�������>���S"OJ��a��)�Pڴ�I�pvY4"O����d�x���T� 7L�4"O���2CJ�K�6��(�+&��ʐ"O�z���$#���WɅ	#j��3"OZQ�t"�&O@|���]:Ωxp"O�)��y�@z�J��Vﶭ��"O�$�@��?EٺB#������W"OĐb�#�#y���s��'tR�"ORUsR[�#�v嘖�A�&���z�"O�h� ��u���R�Bi��:�"O���A���?��ŒK]� `"O0���(&����'���L܍s�"O�8 
�Y��l�,2`
(E"Of��P萴AF�ܳ����]�Ę�"Ol�R�ޒT�@�h�6����T"O �y&�?��b�س`m\�j"O���4��0!��H��ڵ_�,��"O���b�Q��q�w�:'dz���"OrQ3��$���kؓS=�\��"O4$jPFY�JQ5;���X���%"O᩷��B׸dAa�X�s8���u"OA�W@�t �|#%o636�:�"O���$j���x]�Tn�+'x�Z�"O@L�eJ4pTXҡ�&}�4��v"OV���5#-��cԗ..�-�"Oʽ��/�d�l����D�eXLj�"ONEs3��ePl�jg�۪�����"O�x��Q�S�a;�C��P�ⱃ"O.���V�:��d`\L&����"O4HXsl�+!U>q�r���5�.7"O�8���O"N��EJ�->T]�R"O�̻!��W�b�Ƞ��?#�!j�"O��	����4�@�	�%��"O,i��F"�|���O�x�#�"Ob	XF��9R���`H�S�"O|��� ݧ
7�����ٓO=���"O�Y)�ύ�-�(kGd���<�C"O��H���<$j�ī�עf�3�"O.��p�C%\�RDB����XV"�{�"O��a�����Br�Ğ3�.�+"O%�#�+s�0���R�Hmٔ"O�A�FӪc�ƭا.H�!��e�5"O��woA�n���#I��N��1"O �I��ׇ}[� S%�ԚOu���"O� <���QLW�|8��+a��|@f"O�Bt���k:��JJgʠ"O�q0��.� ȩ�H�.s�r��$"O��e�	 D5ܤZ���5:��G"O�I�&gP`�$�7.Y%Kz <��"OrMa����s�Z<E&˪Xju��"O����h���$�^�=gΩ	�"O�@���@�,iI�G�לi)���"Or�{ +�4Q����R��ѹF"Oj�+p&�5xPީx.,`�B=(�"O��j�M�h4 ��
A�Jz�1"O�!	ff�
&���ٱ��t�Ф��"O4�;��׆���B3����p"OΉk1m^[�}��O/�$�F"OִQ��W���q��ʝqu��2"O.q)P/ ^J��w�ʧ3YB�#�"O�I�V%�<G�Њ�-@
�F݂�"Of8#�IO�fLse�J�Vq�� �"O�͢��ǙIŊ��g���2}�$""O�ɛs��L��Eys�H�pg����"O|[%LϫH�d=S�Ƈ7�|�&"O���A��J��D������ �"O��6�J�y��p�gÎԠ4g"O��j K�3�j����;m��;7"O`��`���$�R}8�+U�T��0"O"m1�l@5k2�Yh���V �"O~��f������æ�ȴ��"O����ҙX��  �v�D"O� �q��Be0i�oT\�ݸD"OfpA#�|�J=R��A�YV !Y"O�j���>)���(�.+U�Z�"O��J"6Z�|����Ie����"O��D��ug�%z�M�>�Vy��"O5ȁ�+a� xs._��jIۢ"Ob�8�R�ВA�핡(},t[�"O<(�K!����TM�1N	*�"OJm �`�"i��ܫ�I�#�f��"O41:֊��'oD����?�z���"Oh��"��C�R��N�q�"Ox-�!Fb�m���Pf��t@\�<q�!�\o)���-��
dGM}�<��"���R� Í-F�*".`�<�	�?��jD�b�rl��w�<��P��l�pJF"@�jɡ��QH�<)�Jď�HE�я	�sr��P��[�<��m��q.�0/	�1 !XS�<94�ėn>4<k��V'�1�B�v�<a4� �nϼ�yШN	j�.��N�w�<�g�ئXDҰ"󇏐)�|�5a[�<q`\�@�D�*�c�5'3���!�U�<�!,|n���
��on��c��Q�<q$�v���ڃd�
�������X�<����-�u�BH�t]�El�<a�c�"݋#��T��jS
�l�<�֦�Z�`�����W�D ��DPi�<����i�b�s�A�N�X�#4"�g�<���s��טB���{#�g�<�� �6B'����V�D����^�<�
LHvhx�V$B3�<���S�<�pi�p ��s��A�7?N�S0��T�<G䌈?��j���C똭���S�<AR��uV0;g,��ZHJF�<qB��r�X����`z�`4bJ�<I�kOl��A6(��c*D@�	\�<� �#6ꆧs@�h��KK�68�a�"Of�ʰ����A� W���X��"O����%	;�y�@�ې�d1�"O"�V�� ��M)C���S�j��"O"�JW�����4ף4�d`e"O���5�O01b.T��cQ!	�\�W"O�h��*%���ӡW�=Ϟ}k "Op����^(s��˃n�Gi
�R"O��vK�?}�p��L�0cF	�F"O�0��ك/��Mj����Kc� a�"O^�h����=l4Wa/4Ot��2"O�P���g�Ȫ��֠79ft�"Oz-��J��G�r5-�>	|��"O���B��8۴e[�̞Q��1`v"O��B��LȌA�	��T��y��"O��z�c�E-<l)t��B�$�"O�͛=_a�9�rk�Hr$��"O�u��H
<V*�[!*ɜ1Vs7"OF�ŊTx�������-�ڄy�'��$���A85��{2�H�x�pz�'odE��gGT�r�H���m!X��'�h�{�
�;D�	�1AJ/i ��'ID��s�@-V���`�<6϶�X�'pް b ��vڒ\�g�_�
��'���b��2$u���엟M���
�'�bX�._;6DгvbޘO�<��
�'������)B|+G� @�BLy
�'�� !��
,�F�Z*�
�2
�'q��:���\e��	�"�$p`
�' �5�7�:/-��eݫc|�ո	�'�V�×-�$����;���KK�<�Ui�?5@�!��8�|�2'�H�<ɲ���D�����R�B�C�E�<A@��2.���B�yI����i�\�<��E_Ba1E�/SST��V�<Q�� ���XǯBT?l�zE�WO�<��T�&ք|��
�m� T���J�<��8I!ܵ�a��/K5
��Z]�<��@)g��q���V?Dd��S`Y�<YEb��i�P��geޑJq4����EW�<Y�b�$_L �Юǲ.�� #��}�<9d�D51�,q@m
.o 9D��x�<y��ޣS�FE;��|z�q�GI�<Q�C�.Р���Q�q�E+�E�<ѳ�_:h�����"7h8*�%�w�<�1g̝~qh��f^� ���9W� p�<�gO9V���b���*������w�<�֯م7�B�s1�õr��M!գ�z�<1�M��<%�AbX5zN
A	��v�<�7��;^��c���5P���r�<�c�\/g�@𷁃�J�NQ0��r�<�����CIP�@)=�4�Cm�<I�+$�\q�����E�6�K�-�R�<�TQʜY�̟.7U-)CAj�<�!�
d�,�څlϓnX�� ��Ai�<Y獃[�m0p/˫}/p�Q�_g�<����:`E܌���+T� Ҏ^g�<��g�5;��aF��jC��\�<�fLC�������aܸ��@Q�<d]=�|�c��w�1SeGM�<�&eЉI9�|r2�M<7;���!JT@�<��D�c��U�^��ԦGy�<����qxV�2rJ�c��I�<ip��u���x�R9���7��A�<� F��F���+�lP0��;	�h��"O��j�n�
��# h��s���@A"O�@�$�yI���bGGe�L��"ON�`���0@�[�ݹL���"O���TE�T0pf_e2h��"O��v�5Ovp��E�!W {�"OZو.ںm���:�Jŀh�j�R�"O��IG���`z��aD	��E��h�A"OB�@ׁJ�m�4�K ��
�Li�"O�k`n�S,TiS���4*_P��#"O�	B�D�dF��CO
����"�"O9P�dКw��Iюݱ�"O�H�WHŸ�DJ�+Ѝ"P
���"O~p��cݴ f��34���δ�"O��A���
Fe�d3�\�Bh�iC�"O^!����"L�S��.=n�sW"O�%�䈖�-� ����@�6"OD��%ĝs֨��Զ��8"Oer@�2w���G �Ҷ0 �"O�Ꮡ�H.A��i[�h���ۥ"O����l^'P��˗�� eo�l�"O�0���`����oW\P`A�"ON��l!\�L1��L	:�y(6"Om(���b?�!V�Ѝ,$y�"OP�Rr���5g �"�DZ�R�2b"Oj��!��
Y�+T�ٗ2��k4"O����X�{d�+#�׍]���;u"O\���σ$I ��i֊�1�~܊�"O J��G�Sh�!����&�t�I�"O(A��$8�!�0�G$�(ݚB"Oh����CDy8��0k��R�"O84�D��$��ҡ�6��X��"O���k7^�2xJǠJ�iu����"Or�R���4#��\sq�~�5Ns!�d-��%�0	��{��|�dB?!� �	ǃ.[�\��R�X;%�!�d�-p���*�	C��@2��?c!���>iij��$l� Ka!��7(�j��vfĿS�ν�4 $?!��n첉�拟�nh9�h��!�D�m6X�U�BV�V]���غ�!�uƾ��+�sb� ����!�
�mh�թ�e� Q��A�f͖Y�!�$
��ȋ'͂$��T�&@�,0�!�D�#E�Y�$���\��e�#�͕P�!���r��ߤ6l��	u�Ϙe�!�^2-��@�!+�IW�	S�O��q !�d�Q�d|���?��5�^�!C!��ߝ�>�*Ӭ���2ДmҘ>,!򄌑5+V@��D�U;<8Ы\��!���*��qb�,99�����T"O!��V��}c ͝M!&��iMm9!��u��E;v�2`�{��Ơs
!�dK>\���C �N�g���CJ� �!�94V���%RL���B�D!��)$�B����!bA�t#���0e%!��P!%����&�&FE� r�&�!�D_4�l�j8��M`F�Ҧ�!�dH�W"�(���W9�Z3��N�"�!�$�!D, 2lKqP@X��\T�!��̽i�i�B,Im�@�,F
um!�����NF�,iJ��B,J4�!�d�
4��1�����Z	�R�Z�j!����̝�qF�<[S�	�BON�\�!�� ��N��M�;â��Tu�'"O~���'�8	����BY,��"O�mA JK��&�#����V�f�Q�"O�	vOE�Xe��1;ך�)�"OJ�
�`P����	�3�:)��"O�ٓ���PAj�ruI}�\4��"O��k��\�1�������%�t"Ob�U�S~���W �h�����"O��PfbK/8�x�%��9����"O�S��8���ć+���p"O�cl2'�Ո�ܪ^�`��"OZ����Z`�ҤK�{~r�
F"OT�#��D5ot\أ��5N��p�"O.�@$��1�pݰp&�6C%�r�"Oj)�jJ-��iJ��жb
��R"O^1P�Q�	!,c�&�I ��9#"OĨB��S�tL�$��-�Ҥ)�"Otu��ژ�BP ���0b���xA"O���@&�f�*Ah"+Ґ{�V`��"O�)R�A�NK�]Z�i/U�8�"O2�cw�P�gb�rfi	"T:��u"O:��� 
:�`�Ҡ%S?WM���"OVEz�a^s�����)�"UK�"Oꬃra0iq����M�T��D'"Ov�K��� �r��2��$:�!�W"O���KQ,=��i��]�(9FXJ�"O5a��F�f�>�����;G.�l@3"O4�E�?(N� 
��v��8�"OF�C�!B�K���k��H3�$��"O��L�<�����	$(=F�ط"Oj8�JO4x��F�۶z&0�Ȁ"OmI����Z�^=�RMF�"O��N�2�(�g�ڇ�P�P"O
h�1���b��ۖu�B�c�"OZ4�F�	b�"�*Z(9w4�b"O�u�1�
.��Ui�iW�uJ�:&"O��g���ހ0�ciQ&f�u�5"O�b�To��#��K'��8H�"O��A��8ʄ!*Ë3ꖝ�"Of�F�$��l)D��O��x "O �[U�F�Z���$]�Tz��""O���m�C�D�� �4uŜ4�"Ov�(��8��0���^�:d�'"Oऐe�-��URu&ґx5�2p"O�m����>Aaf�2P���q"O�.ќ[�F���"z��3�"O�"v�eW�����>5"��"O��zǅ$1Fh��A�y�N��v"OL�^�3�8�1d�F�\����"O���L�dxST�>h��i�"O��	A��+��%��
ܾq����w"O���$��)�jk�'[��<Ba"Od�E��=x�|�&H�/i�J�c"Oִ���TYqF\�F��X�"O�Q��Z^~���Y�V�l)Q"O�$
���,|0���E�UP�"Or@01����S���Xi��r�"O�H�e��R�HųcD�kkd��"Of����@�Ru�X*��ҩ}a0�"O@�q�
��_����h���`�"O&����3i	�A)�!����C"OTe�5	�6�<��&ҫ=�
嫕"O�4��K�.��&��q��5��"O����P���L�E� ��=�#"O� NE�&�΁7R0�q��?�b�hF"O�@�e�:��!���g�~�"Oj�w��+9��%���	�Х��"O0����	�%�"(8�NE�]ͦ�:�"O<ܺ�̅�8��]	R.Y0��*&"O�$�eO�Z&y��.��YW�q��"O���Z�~t������[��bq"O�[�*&$�~��A�A2ap"Oh� ��?h{D`�nY��ؐ��"OX�.':��`�.6�lD�E"O\��AK(�$*�fɧ<��R�"Otɣ�e�[p<����ͺ��"Otw���!Ȗ�Kq�(v� ���"O:���\�825 vLy�Z��"OV�2$-P�A����]+l@�cW"O ��fj�0���VH�n��`�"Oƌ����Sm�9��Y�y�Q#�"O��
ޠL��(�J/+gxi��"O�)*"(
�B�$���f՞���q"ORyxG��,P�8�)�˖�>;""O����`��s���ӫΤȀ��"O���'^0l $�R됿oJ�r"OȨh�	�0tHI)p��(4!l��"O�	�I��R�� ��y���"O��g���C{�X:qJ�x�$T�@"O,� �U�ndsvh0`���B"O��+VC� ���� �@��,�s�"O\$�E��R�<�G�=L�u��"OԃbM�	�D��&^2�$Q"OT,�A��E�t�dW�r
jii�"O�mY��۩dn�ʆ%�	T�\Y�"O� �	�e���Iwf4��P�r"OH-8�AV<V�@3�ͽ,�z* "O갈�����̫R
��/߄�q�"O��c�K�j ��W�
�p}��"O\�bLC&\����U`s�q�w"O�)�Rߺ�{��Qe�\��"O2]��$Q�f���̮����"O��U�>�  ����B���"O�1,�oΡ�"EN8B��
d"O��$�U�]�1r��gZ�7"O.}�qHT;zG<l �T�=`�H�F"OB����c2 %��$ѴzN��"O����I^�*ԠI�&��Aت��q"O��ె��G�H�`��F'^����"O6ĂF��6�в�l[���8
&"O|yZ`ꏱ=��Q�k�,�\�`�"OT!��oܦ>�H���\�8��d"O��B�i&zq�E P�jĠd"OVl��
Ͽ(h�Y7בW�Q6"O�yR�M
��Ї�D�bgl��"O�PC���+(�Z��E!fd��v"OT�ڕiC� ��y+� ��z&|x"O �I�Ĕ�<��K`S	
y��"O`�2�瞽PUԭO���*�Ѧ"O\)���ڮ;o�	�%D��0�e"Ox�J�.�yKFc7|�x% �"O��t㙀xw>AZ��[\I���"OFHH�� :>*)�����HB쵑G"O�9"�G�������%!6bEB�"O�0��@X!,y�ۇF۟kSF���"O.O(t "D���#8(l�p"Oڽ(SH����y�zXE�"Ob8��Es}��c��^�v����&"O� �-���\�#rp9��xh
��6"O�4����)~n`��p�:q��UT"O6,p��<m`a3/�D�P⦀��6��#�'0FH(�a�fecw����(9
�'U2@�u�1H�N�*�n^	Y5�8	�'�0���˒�V�,R��%�X���'���r��F�{�$�6 ��c!Ɣ:�'�|�Rd��u&�ʰe� �'����c	�}�*�[�*�Yu~X��'������@� 4�m �O{�|�'j�;f�K�q�2%Ac/�*�N��'�<)Q$�SS��,(�"�	�f$�'!��B�<	��c#Ǌ����	�'J�����6�$P	� �^���'�>�J�(ûm��H�E���d��
�'��M���XWBp	a�	�Zo�
�'��P�	��L� ��^b��j�'ؖ�y&�':���С�J=�')d���Dխ[��%��V�|A��'�Tp��풉[0bl��E�~�c�'Զ�3IC��*����:h#�a;�'���ޛ?��4��e��g��c�'�����M��qr���Mڿg�U��'�f�a�j-J?~��'���M�z��'٪� Θ�:��	1�K��;��$k�'݆���hÛw��X!4b;�D@M>)$"�;�@�<�}Z�`�5DJ�Z�-H6g����ǌ�e�<��&�";����QCM
?���PM�:kT%&�T�!��������)�g��!�a���8�H���y���Br�O�	x�+&�Úx��"��/'������x����JּY�Z��oAy��1��.O���
��|��;��h}�(˒r�(��M-%�A��'���y���:1�8��	${<�Fm]���$T&"v�̹��Z�qښ���S�� �`E�N��<dJb��"�@B��.6���r	V�}�@�oIi�F�2�ϯ(���̴S��l�%����-Lw��:�O,kWRpq�T�:�}b�Խ8����GJ(��3����	��Q���.G\��P��W�y��x>��J5*�K8�Lz2ORy�uEz���<ot�*��@�P8	��j��>��	O�o������-�l�#��RF!��.0�����]<�����{ܘ��@C�?j4��ա*86���M�/�H�׍�R�4�k����t��G8�y��2xz�0�2����|A5f�D����狂/��C���Ph�L0�Ox� Dy���F�����HF��7�ٖ��=���8x�I�Њ
pd��)A#C��1!#�`P�Z���~�
D��s8��P/�&O��@����<H>�LX��;����]b��H�J��r)B��n���N�?}��iI9:d�����![؀��+6D��9�!L]n��@M���MI�E��?�8��bk̂���JbTVL�3,#�'�y'/K3`^�E
�eчa�B]��C��y�g�,l��|ar��ؼq. h�U]�Xd1�pa�u+f(�����𡰆�a"�j� �
<�zr�G��
X�dÌ ^�Z4JE,�!�c��-br����B�JH����>�<��d�Nyniy�/�a@�(y� �"�qO��I�G����H���
z��4{�$��~i��L�e�c��]��`�0�R�S9�H���Pߖ��/�+Q�aK4��q�>Hj%����܁j���5B:����"�Sj�����LuY�`�T=j�R�m��3�!�Vj}4!V�Ւ.�ɠ���rxq��gS�e�B�@ݏl��eCg�h{:I��H�y�,��#�
dg�ap��Q�z��Y�yʈ�u�$z���cN9E��5�Gj�9X��+#ǄO3��꛲{�����9(P�6���]���TkZ5�qO�]�E�N�^rr����5t��f��Y�����[\��oD:��ڴ���A�ȓ#�l�E"
b:l���o�D8�� 2�G"Z/�x×[��Mq�"��rx��w��<��%����Qc�\�$Kx�	�'	���3�]#4�\�C2���+�ʨ9��<�9��P�D'��W�[hc؄K�G��hOr!�̑�Z�8��xQ�ɛ��'`|�p�
�z���z��9� �UZ�J��gCة2��_)?7f�K�LZ���a�'���QC�(a����լ�+dZ.ݩ��,�$9���C���S�,U�������^�d����\�j��ԦW&$ C�	�aD��∕8cpBQKaR84�V��,�P�+6g4?E��'z�)�K�F��t��U ��
�'�����^�	;Ԅ�4Q0���'�ʘ�RX�'����͋^�|��*S�m����)[�q�!��85��Sa���B��ţ'.��7�!�d�����g��5lت)[coD/Vh!�D���`hX���	��h�ᓾ5\!�dT!<�F(3�@ 8��	{��רlI!�xs�谕KO�,�P��f��V�`B��7����D�@a[��(TB䉽H4�P']+P�0�i ˜)XB��-P�4�Cj
�T �f�QP0B�I�M<l�*�ŗ�,��׷rB䉖\��}+�m��AFI��.ɷi4B�	2m�����ПK&`rq
/.�^B�ɿg�|��+.a~��R�IW�'��C�	�9��1೯T=m����W71^�C��|܀4��Մ4ʹ�XbgX&�hC��$/��!���4p��]�&
YqnC��n��j��:q�b	��GR<D�4C�ɍ�\B�D�0,����KE�t�,C��"5�-��E�(&�@��;l�C�I�*��aG�P�E���Yr��!M�B��3A��Q�H�!)������Ɍ<��B�I�|��BVoޥ�M �Α�k�]�ȓ
Y��AE�K�"��',���FQ�+�k�b�b��@ߨz~�ȓ$���R ˈ_ِ��vɤ%�e�ȓ_�\Wa�9�z���G�-8�\��0�V�R�GU�e}�XBv�(Il��	z��tH��T�9*g��^����ȓ<o-�q)��x�Q��#	�`
؆���zv��M���RB���D:r�cN>Y
�b��%�`@;�z�е�HuɆ�	�<��,D���`�>��Y�0@Qo�<�w ԍ.6~�q2�@w������W�'5?%�7�-e����c�;I\��U�'D�<�`V%]��xdꓣ��tz5d�<���eц5:ĥ�5@%�p�Ňċi�B䉭9;(�y����� �C��$��O�����q���f^RU�e`��vY!���.�r'�G��C��<\!�أH
��`�K�-%�Q�b7#!��}��4���E�c vy+�c!�d�hm �'Tl_�(�$��D!��:I0l�ȇ�;ݎ5�(�-�!��ʰ=�L�s���'����E%^�!�V#,F,���X�3�VY���^�!�$D."�iG�1���8�N8Yz!�$�.Uq@���R7�~(���T!���k���Ӓʕ�4���
�@YQ!��yA~ԙ����0�D)FE!�\"*������]�KdpH��R!�O����E�B�7����.#J!�dƿ/겑WmI�%���a2 !�$
eX@5�0ѹ[��%Kt�@ I$!��60IAI-h��	�DL�<'!��q����g�=E�Rqu�0�!�d=[�P9@�R*i�Q$J�6yW!�d�K��YI�G��EF4D���4d!�$�
`>�M:4�7!$�IAƎ@!�� h,��n�� ��i����4��X�"OayҢ�02�� W㐙W�|=3�"O �sff�`�h�8�(��Lpu/��gg�%�=����Ob���5-	dh$쇨S$\�H�"Ob�떉�xҸ}� a�%(^(��-��o��d��[�a|�Ѱn�L%��ݏ�h�b����<����x��Z�]x7� 6w� �a,"8Lp(y���V�!�$�c��;�+�0V̨z�D?3ˉ'a��I� ə|c�q �Q�q&Q>y�	���U�A)� Lb�l�5i(D����74��Ba���U?z0b�e� i+>`s��ެ��"d\zb?OxlANӥ~����.v��:A
O4�8�HV��Rh�q�<�^�[�i�%�n�Aq*��O^ы��9�0=�b�K/���I�`E&LH���SI8�|�ׇ�"	�֏N�O#�����'��1�/͍��@�Џ	�*!��+C����T:0��"ՎۺO��I�uc=�]���TH�)G���貫4�S�P ۧE��*I��-c��B�I�v����ՙ!���1&��&L�8����l�N�1���b��i)R�)��_��/h
diŇ�]��T)2cY*BB���in���T�2KI�>���	]�<�y �D�/���ë�qx��[	@?��q������x��0OX��� ��I���Gl�8��9�4`���JE	`������!
��!��B�ɜC�.�J�f�)L�傠ՠ.I��S�>9�ڨGP����ߧ[��`9����$K �����?o|��ԩ֦�y�aPzN�T�&��b;�YLX���"i8�[��mA���Q^p�|�I>b@X+e����	�2 Qa0GZE<B Ho��1Nզw#�����Q�j಄�Yv�BA*�b�-,���y�|}R�*C"Y�,ѕ���~>r܄�	+�nQ83d� *`����޺^�,�!��[�@�>́VB�'8E���"O�E� ��q����!a�48
}Hd�>)�#¯'n~4��E0kP
�	5�'�`ň'���h�=1�������h�L=y@팋g��SA������)��Ĩ�Af�O�-H���^�g�	�V��7��0Y���w�R ӰB�2�
ś.$͔Q��Ե	H��#�,T��j���:lNY���`� ��p�݈Xt�H�1��g��ĝ�Yw�X�qߍdy	޴n�|\8�&��,AI���4������ �$
/E�`���F�� ��=aRc�}�X5 !�YD���
'u���늆J�����V�,�+"��8��QxU�Ƹ��%j��R<"#qO�}�#q�E�QP�}�,�'�F��ͅ�x����$�.L(t"��F��\�ȓ���@6M�Z�.���/:�����3&Xr �ׄ3��l#��P����E��Y$ԖxH�r� `�^1�ȓW4��feE�:r���q�$��ȓg`�L�D���'|�8��ō1H�\�ȓd!��u(+'I�Y��I�J@%�ȓ|���('@��P�bir��Ŏ(�zm�ȓu�ԋ���3
%��G��|x@h�ȓ �(8Cq�K�"��@H�cJ"dS\��ȓm�@]"%�Z" ���A� O�PFd�ȓ	�*��� O�F ��+U`��؄ȓ��ّ'%�='Z&(�ge
2g� �ȓG8�`���jh�����9k��D��3\z	1T	]=V�t)���"�r0��o�a�f�1
״�x�I�5�I��E�AC��T"x�~��v�K�Fä���Iy<ա7j�~�+�,�Z�"O�Uq���k&pЃ�9P���"O�,;��XjE��O��P��"O��dĊ?�Xy� c��R�"O��y�$#d��́r
*	��2A"O����#��ib��#M�V� B"O�0��l�")a����ԦG�ܰ��"O�h��JX��DP�Ɗo�t��w"O� ��3N�� (B��.��	�3"Ob��!�F���3�$V	q��}��"O��:�HS>Ov���B��6��@{A"O�f�èq*U��"Iab6"O��B��D�e����i,P�I�"O~IqQ)�h�����
r��"O��F��k�!�W�AV#�S�"O��0'�8۞ �U�\c"O��Ɍ�$*"�Ҕ�(t��8e"ObQ�ƀ�0Al,��U��Nm0"O\�9�
�?I�X=p$�<%�,�a�"O�!�BK�< �y����t��w"O�i+�N8v��a��(�+JF���"O�<���>?�$I���ų�8�"O&�+� ��z��J��;F�fȸ!"O�2��E�����IѦ(� P�"O�C+H�]�(�;ʂ,�"OR�p�-y�d񐗍H;x^|Q��"O��14��r�
�sBlL9.2���"O>$J��*Kx&���+B,'�l�U"O��y��l{��4
Cw���6"O�9�#�֛w�M�6-� Fm.C�"Ol�9P��8.� SL	�T�,r"O:e�#n�1y�✋��]�*���"OxA�a�C���
�%��^h�r"O�gF_���w���u"!Pu"O�L��&�7����Q�E:qT��"O�UЁ!�T֮�`��? mJ49�"O��a�/C�7�L�
�� z�J�p"OB�:!��(W�"���Nݣo�iY�|�n]�n�mQ�y���aȚRm@e��Dެ<��0L���y��0�-0��\
0�p�n��4���K<�BO�%m���'����׹ay�9��M
�s�8�	�'��\�e�%��!8Dhϗ4�8P�lS�Y rI`�߂��>�' d�HQ�r�ָ#eFy(��CO�(�JB ��SJ����J)�X�b�w�p�rC��	=�!��ɸC���Z����p���2���s?\B�� �4�8Z�0�M�M�d ��\���rV5.C��>��0;g-H&
r�����t$���!O2r����9����b+��$Ԉ2)D�8 	�.2A�h��N�}�+��LJ��8?.nA��j	$J!�x�� @Ȇ��3b���P��7�<�nIS�ܰfdJ�uI�EFz�MR�pp2ǄI+PaF<k�EK�&���"��\�3v����%�!���8� ��4k�� ��Q�Ƶ�p��S���L�
03� ��0zps�χ��H�'J�:MtȺ�ֱ/�<l�����y""�*p�<�q�f[�!��k�*�e/D�:g(�m�y"b@�>r���!�O�:�EyR̀�^:�����ݜ$���ȥ�@��=A���_� ����Zv��@���e:y�#� P=���	��P0&G8����`�&��2�J�cڞ��T�(���|��8q�# �&+Z�õ@T�=ͦ�>Og���+C�tp�-��RͲu�wl!� �B0t$��#G/0T$`q�E�q�<4+�b	�t��5;��Ôs[p2���kޡ���X ?{�9b䞟7Y�t�&D�LP,�y堈:�\�>s����ǈ�@�ڡ�.K*u���獊=t�֝0un�Gy��͆C�n�S�H�nD�%���>�p=!�*��f�dmV/S�1���#Z4DH1𡕁s@8tb�*��i2�qD�|J��XG���eN*1=z0������'<�YU���B"O��(|L��a��\4��o84d)��ڇZ�122a��Ud$C�ɍ|���!��<n�d	�ʝX1���i��d~��KƉ'����O�~���d�țw���j��ؓR�t���[�l��
�'������I����v���c�P[�)^~
���Lh�Q�!L6s����w!@K�'*�$�RLU���SfHHYZ>Q�ד2ŘZ"�WH[���"��t�-���B�T�ta��%N�t���w\�" S�'�^��ċ��n��0Z.�6�p�؍{�I��x1Xܢ&$X'.P۷�� t�"���ä?Q�Z�Dɻ���?@b��W�4D�� <�yA+Z�6��lB������E(C����3��J$@x�}� kI\�:��2�+pޅ�	D>wh P��eIwni��0D�p��ey<j�!�|�[-�6z_q���#2lp W��q���W�'���a��[�� �W��_�����e�b����Z}�i��M-1���7�/�pd�d�.1k��bP㞌~aa~"nR7}<a%T�59��!�	�	��'�>��\�!h�l�Fʨ'iv4�K?����=*�!a�
X�.]���ybA
�X/jm�iԛ%�ԍ󤃙�$�\��"և3�@�I�O?�IS����/�/�>�	Ƃ�p��B�	2��c�(Z7>t���v�j�I�p�D٪��K��p=��+�.i�x{ DO�#+�]�f��w�<���K���7��0A_� ��&�q�<Qe"��Ri2�y`�C�b^��c-CZ�<Q��P:7H1 #�Χ@�^U�C�Z�<IP�S
|�P80�T432��s�bEP�<IS��7*t� DD@�1��pK�QN�<����&��E����1Y�&i!MON�<���5y���2@\F����Cc�O�<�q��}��g%K�_Ex�F�c�<��ŗ9d�ȅ0�nҸ,$�E�X�<�#�	5�(�	�C�x���L�T�<Y�ˈ�eDP��4R��I�dD�<iV Qq��i��
݈XY��3([�<I 	<#�5:�j�2&,"���@�j�<�7h���x��Z*X˜�)u��e�<���T��l�S��*{�<צ�_�<9B�P�}T4�Z>l�FI�@��c�<�o��%���ЬE�H}��f`�<YG�T�LeV٠���}���g(h�<ٱ�5=�HQW�I�So���S�f�<�Q��U�Y�)P)���F��{�<�#I\v�@�� ğ�6Y��)3GN}�<�/U�:��Y�4�ڹC^ �$z�<����SS����H-ᕉ�c�<��Ju�lm�T� PT���E_�<a�Hӟ@��A�ǁa��83�_Z�<�@͑�ZnI����9��`@P�y�<I�FQ�M�0�K�"��4���	{�<B
T2��3v�M	U-v��� �{�<���@Bq�VH�:.�k7�q�<)a�������#��6�n�{5�WF�<�!\�3�|Pj��0�:�ك�I@�<Y�c�6�� J��_H��Ѷ#�<ybHd�zD���A����+��O]�<���J���v�@1=�R�	�fLZ�<��
6c҆m�OZ�J��0�
T�<q )�!^.�҄̓*k���AV�<�P�O�Q[���#%فl�8�:t�Q�<	BVcp�PU�O�p*j�Z�!�R�<��.I=)��g�?0�NeR��YN�<)��+����@a@�J����v#�c�<�u��>�4���ʁ�`-ji8��NP�<���1!&�k��E3o��ԥ�F�<�3��y�6�q2��5L��)UNG�<a"LֹQr(@��O\��y�MRG�<E�b��@�G�W� �pծk�<�G�	�N<�%BS��yG
�\�<��n�u���� �֌ PѫHf�<�'��uOLE4�C�bRtZ�#�b�<�S�G��6 )�jx}hPX6��A�<)��V�m���Q�
fr�ID#�B�<��D
�(��E[�DK�,�dx���A|�<!6�2n]Y�i�2 ��r�{�<��.ҷ�*��`A.Bդݰ����<� Leꐠ_�`��C��S�����"O�d��_
c)� ��H͌[����"O�dYF�¹.�<�� @�]����A"O�ID �2慲q/�%iw�Ő0"O��kC�p7#C�P�q� )!�Ȓ��6K_5E|��c��H	!�䀲W�´+��O1,�4,�e�!�D��mFT�r�$M܆M@�N[� �!�۴?�i�7�7/@����.!�>l&�X�3@�pg�ݣh!��M9Qf��A�L>��Ԃ4
Ĝ;�!�D�zj��#�nZQ�eɥ鐁;7!��S$LЅK���	��XY&'��f*!�D̙g���Q��
e�X����T�J*!�D^	3�u�R ҙe�f��M<g!���H�NԘ��z�g�&�!�.;�	p��S�D,�I��!��<`��Y2Ʃ�x���:�5	!�d�|�|�!��	)4	��S +�!�F�B�l��cӾ]�P�yS�Ŵo�!�=EĀ�����Xr,\;�lC-D!���:~̠u��-tb�푲aA�!���6�T0�IETv����.�!򤛮fe �4ϛmBE{�5�!�dN�$� ��7�`6�Z�A?>�!�D�ܙ��Ǒq���g�=�!��ɤ$�0����,R,�AB��(=�!�DD1B���� L�4�3kT z!�$������.˧>�3#���1!�Ě�n'�����L3?.Q�1Ɖ4&�!�d�4�%ʳv Kå�y!�E� g�D! �,t(`�J^&i!�䉨I5�``�*çv�"�:�
T�lV!��U��4ѐ-\aX�JgI�(jN!�X�'�e��iܓ?t��.�v-!��L&�t���P:�d�ʑ�عi	!�d�(=f��+�6,����g�D�q�!�$��pb��B̾CZ�`�����3�!�䂖W ��q�H�'�:����'�!�$Ć�x%����b��tsGR58�!�~ lh��Պ[1nih��{!��!Rh�V�֩�&Z'�E�({!���
b0t	���cI��;^�8$S
�'	@���H$4
裠�B�`���Y
�'�������2,�iA�Em��S	�'�yYoW�=ݼ�!��ɞ5P���'-�T2E���1��� O�6D~���'�Ģ.֏yʲ-s��ӊ^\:h��'��r����T�lM�Q��3L�~���'Z6M!����yT �
!�B�(=�'�2d��&E&x�@ ���(,B��
�'Y�MCj.	�CK�/�@y�'��"�dٸ�xh
�Hґ_��R�'E�y�t��W�(�Qɏ�a��t�']����d	o�^Q����(Y����'M�p��� �~� �R��a��'������
?ل{�3YqzE��'���@�&vo��B�C�5mQ8A��'/b-�"��D�1Q�L
�a��Th�'�
e%M8Mo@�Q�GC�	-�K	�'�X�8.H�j <`3�"7&�-k�'��$���&��8����(D�qK
�'-:Q����3���"+Y5t�.j�'�������.Y� 7,X�k�L�*��� �H��+JQ�%!��X�ʀ1�"O��kv�,0
i8�)�n�<k�"O��j��
� ^� ��V�@���ض"O�Щt�"������4�\���"O� �@�.�����	@���d"O� �Aɔ��$=s���>��b"O^���l�B�ZAH����v�H��F"O���e�:1�( z�i<L��0W"O��V�R:�J���)�z��|z�"O���	�'.4�鲇P��d�[3"Oz�i�E�k�h���*��SF�!�D�֛�Pz��,���|��f8Ɇ�z�͍�9����/3 ¤�%���O� æ���I��]��m�3�R$V��m��Q� �����o���S�O�:��g�֨�쵉 �h	 ���~�h�b��c�ҧ�����	�;1��Z�a:Z��	P��^p�Ա*�>�U�EQ)TS �s�C.k�Ԅ�Մ5Z��\�h���sӐ �ܯE^"i��lXP�؀�xR*��a��O��\MBf ��IkHxش��FL�I�X�HRS�#��|Ҍ{�d�J�������3:>(���֬�?��k�����-Y�?1��0��)�%Hŝ���y�(ς+���8}�J�?��S2_�8���9>>�(ѕ��S��p)�U����d�Ob�����|:��?�"�s�A�9���L�%B���V��a��}�]*��:�u���ghG<N,<�;#��$Olrt�G'�
x�t�����?33�M�Զ�0|B�ዞ[���?L
L�;���	 >�\�{Ѵi �m{��)�(�KC�|,�lB�%X�udЕ���>iGsӀ1RW&)a�a����{��d ��ΓLj=h����y2j�|�q��	-�r��|����%��<s�A�*� za����$�4U1 $�>E��
s�՚�	�%P�����H��y"'-y��㟢}ڰ&�-u�&�T.�H.��a&���!���9�S�O!X�Qn��sq(D����g�0a�5&��(�yW�Qr�/��@ua�1M&��>�ulS�����O,��UB�� o&��V' �P:G�xB���O��pMXЧ�/�~��ŏZWV�9[�����'�lI��V�ul��Q��R�r�N�S�'�h�U	ǯ�L1�G�eg�H��'\r �Z����jR?Z�,�	�'x�e�0�� Rh�@r�֝R�Qp�'|����q�bD�V�XQ��'���@�زo@$!d� �b�d��'�8��L�h0Ɉ�)a��H��'Į99��� �>p�p�0 R�H�'Xd
�;�b�`�O[�M��'�C��!G#�ifG�P�~�R�'p���CQd��L�OK�-�'�0 �%��
�ʬ۴�	�F`����'���aQ�J��A�A��nC���'eF���k_�����AG�*P��=��':�P�BD��P��s��|��'����ށ �TY��/��y">���'���Y@ȠM�}�2a�!�DA@�'���s�g0�,�aa܀E �	�'9H F��֢�*d�9����'m�т�����w���GHH��yrJ��5jCʑ6$0��GȊ>�y2�ů	�p(�����E��Y#J���y�b�e}�vk�'0��P�5"�2�y�J�v2\�f��ug�)�����yB�ۨ Q�B\�j��ؐ���yb`�7܉�f� _�b4�e.��y��l���peŮFqJ��j�:�y":E��:$ƏH�X��Z'�y��O�c�`}��OAf(We��y��	"�h]+#䅫ܢ���h�R�<Q�)(i��i��6RL��xCd�<� P��ţJ4n\4�0̢ ���"O�I`�J`���)B|�\�Q�"OV�B��J8P�$=9D@P����"O��r���n�3�!;Y��4"O�\z��ݠ4��1ʐ����`"O������7Fh ��G�M-����"Op�۠�!4��	�F��D����"O��� l2L���CEE'���"Od����C�cv��QN�m=b�" "O�m�&Dq0�%�D(��+��IB"Od|�p�3;q,X�X

$�R�"OxA�+��F���k��(��ȁ"O��#�ˊ�`����!!�h��"O���Q��{k��ے�x��i+"O�ٕ!λ`�2 ȗq�@ErC"O�H�7(5Zܘ�%�	���q0"O&�bUhH��tx3�@}9�HK"O|c�h���ʓB�7'���r"O�y�#`�3,e�Q��Q�"$IG"O����o�w{ZP��Z�Vl��"Ol1�d,�
�8b�P<�Н��"Ob�r��
�Q	���p�xI��"O���5���J �	ڷgژ]v*��v"OqB�M�)c�C0^��� D"OZ���,�?Y��uG�ƻHj^|�6"O`�ӎB�Z!T	���\;I���C "O��]3tgŔ"#��v"OĜ�W��~�Z0L�-7}�q�"O����4i���O�p9�4"O☈�`��0n��H�L��ܒ�"O&�A��{�d��v��r	:��"O����mҩF��!Ʃ�4,��I�6"O�<A���CH����ovrp��"O&�34g\�Z�pLZtiI� ���3B"O�=
 H\�m�Z�:Ӈ0i�4�#e"O���QeP5d��%HV�ԅ��d�e"Oh�.ϭ�r��T��*�,x��"OPQ���	�t�0��K)Uu0���"OHp�ug";�-����,��q�"O��c"�("=P| �
��p�"Oؽ�ƨ%4�]���^�K�R��"O���(P���T:gL�"O��#�3/Ȥ���@O'L�~�BB"O�a�ۃ�N��쓛H���"O����b�<E� ���``�"O<<�cO� @z��kcK�-k�H�p"O�J2��$�X�9B��1�A�"Oް±L�&p1���:0z](�"O X3ƌ�:��`Е�֝(1 !�"O���Ճ@z*�����f'Z-X�"O,���Eq�<��ɼ(�a�"O�{�eB�o_�����T�=t>�"OցA��0%���1Ѳ�2E"OLhH�o�|w�h�d�����"O��1풠9���������cT"O��zS��y��X��N]�Z~�k�"O*M*ϑ�ۚ�;dLZÒ`�"O];d�A�C��1�.[�)�5"Ot(�&
��{F�
b��Yɗ"OVE8b�S�[$=�bJ��2z ��"O���u�F�]Q�����B�ys&= �"O 0�/���t������P*WHB�I�c5#u�R�c� 1pa�L�{��C�	�(9J�+=B��ce :b(�B�)� (��3�Ӵ	$H����"Oވ�t�&*�q���,B~��W"O�T[ oڼ"I���GIG3�u
�"O�4Z��`Ȩ�[�癅c Tӣ"O^Mi�Ǘ�)� �+�&4>����@"O�\�Q��9E��=#�`��|ר��Q"OiBaO�nߞ$yfo�������"O���\?<'�i2�hߕ
�L�Cu"O��+Y���QM�~�<r�"O��0EҖ4�",����1}���7"O�0�!�qt��a�&^���"O6u�sO�

��u�ޔJ�1R�"OPMx�-K�(3�ř� �]��iCf"O��s$��Z�ȝ�f��g.��"O���ùV�T�IԌ �I�87"O���q(�#	1p`�u钃=:���0"Op��+��QR�8��A�B)��Zf"O��CҨ�g���D2P�I0"OBAs"G�]oHU��-�%
��p�"O�|��⟉9�u��
Ƈ7�XA�B"O|�xe�ϖ(��
�c�ar�"O��ZФk�x�� -޴9D"O�yJ��-(7p@��frҙ8B"OB�P2�	�J��1!˶cp|0��"O�}�po I���3-�3^`��y�/�Lf6��Q���3��t����;�yB��FWr�da�8(kR�ju����y��T�@���6$����*�EM��y�K�p��RT��ga��yHӖF����6n-�reP�a��y�$�<��1��=~���A�y��؍\���X��
z���`s�
��y«��(P�U��o|^\�w��y"o�>}�� c#�&`f|P���0�y�BɵOO����ь'?.$K�j�<�yB
�,Ơ8�ݢ �2uM@�y¬S CE���"��Xv�Jt�»�y��Y�.�[�A��
����@LN��yB�R�,J�c߬}�2�R@�?�y�� 3�!�!o��0�#D9�y"BĹ|_�A�"$�4Y�D{����yBBI�-m�eP��'Q2}��.P��y�_�	�k�Fj��& N��y"B(:r�q�D�>f]��)��y�k�&JL��RJ>���c�-��y2&�#�V���C�#J�|�q����y��  0����D����h���yRn�?��!d�*Qj��J�yB�9]~����@5H�T@�Ņ�y2&�&�8��G��B�R5��<�y�%�T�Le��� <��9SA�)�y�!Bu�0�U-�%*�d�i�����yb@�	WC��@Ԣ�(K��BÍ�>�y"D,ir�"E#� ��B�K�y"
|5��)+[�jE�'&��y� �D�X*`�͘=���UG	�y2.D�]����/.e 2�E�H�yZ�X�	�DԞ_8��+ìH/E��y�ȓOߒ��̔7S�8���I�=1���ȓl_��rU+�8!���
d�X�c/V(�ȓT	@Q!S��AN���U	<1A�T�ȓn�m���Jm����q��/����ȓS��w�H":e���D&,�����&����A�W�D�ذ/߽"TBȆ�S�? .�k*(� �S�(ʜx�l;t"OM(:�h�(Q�:.\�x)&"O4��+��0#�D����eM{�<���L���{Fm��}�5�`�~�<y����BM�Tgة=ց@%A�x�<��߭d�������k᎜ꠦ\~�<�P/@\�{A��?��t�s�y�<�1��x�T�8�.6"�0��_y�<�c'7�F����@5{�j��_�<���ɌsB0b#��`Ll)t�E]�<q/Ƭ-�xL�3�UD���8Ѫ�R�<i��%4����"fNhj�����N�<� K�$�H��Fߜr� 7��L�<i`%͕Z� ��ƅ#��|�G��^�<9��
�#ֈ�(���F���E�]�<��!�j��98�%Y�f��%i���^�<Y� �**Y&��5*J�ة��KE�<��	
8]��)b�1�x x5�A�<�Ǡ��-��y �7�p�%��w�<��(Ǆ� ��Ƣ�5"�]u�q�<a$!ܩ΢��4F�pg�H�<��_�DĒL
c�ї1Dd9A`K�<���� Š �"DD��xӒa�`�<�g&�*O�|�dh�p��V[�<)儋_@�y(� C�<�r4��|�<��W,�³Ժ.RP�4�u�<!��+
Fp���R�^U夀q�<1C@��c��U��H´b��]���o�<�fU�Q	d$��f̰&��X�%�`�<���""�Je���,F����D�W�<�g-R�'z�AE��?20^e# J	I�<����Nʦm�6�:IK2M{���l�<i3N�<��)�_�\����u�-T�\뤭֒"�l��0�Z�r��!�%�7D����)�PlD��j��*|x'6D�h�#GF(*�y+�◬3�4�I �)D����P����6�ִwD�{��&D�d�C�K�Rl��EU�f�.m�1�$D�,�`���sߌ���NƤj��g#D�����
1�L�}��у�"D�d��$   �   [   Ĵ���	��Z�HF	�+:��(3��H��R�
O�ظ2a$?����0�ݴrf�VB˖�	j&� C&�٫ M��lAFq�
HlZ(�?I�')�蹟�nX~2-̷d�^���Ko4�9�ʱ~�<}�I<Y��b���)I>�',��H��8Q�``h^�]��ƬȽ����p��I�3)��^4,�ԃ3٦�h/2��t��4�a�4"Q4wj�0�$i��5G�ʓ'��*�y��հ#%�G~�@Q8 [�Y�S�3�d�c�(`Ḁ4ȍc�8�u"�i �䑎l!�q�$�O���Q��J<�K �՜[�I��_��00��GQ��s�|R-Qo 2�+$�M�d�X�"X��ϓo�>"<	��,�Y!��j�l� K�X�j�)]���f�
q*��R�Q�L�A
S�6�v��ŤK�}-X9R�;}���h�'���=��
�>	��$)��f����Vڦ  �I������o<rP���D�/+�z��� ��C�b�Ѓ���;z/�����C�aw>�����eՠʓF�x"<�� �I��­��	"S$a"VK��B��)ɰ�	
%��(-�?ƅ�<�!��O
V�jD�f�t̓)��#<�6%-�O�r]"	�&�W�#J͛�
~�����O��[I<I�O��d�]�`�& �# ؂e��0�'�"Y����Q���~�硒!|�iY"Rg�E�d
���k�>+|2˓0����`PN�	! ��9�M�1��<��R�� "�*`BŖ�q{Q��G��#4H�d�< �2pc0j<YC�I�� �  ��ı{� �  ��A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�ou�!Dy�'�:� Ή�B�\O�|�����<a��$�+q��@rsI�E�f�W�]�1O���$���R�W����FޜO��'*(#=�O��)1�h�Z��K�`)����:o�.�<�J����<4���y`���`KR5��O��Dzr��`S��o[X�JC �+�lԛ�#D���5�^;Ki�e:	�L�� 3 �6D��@C�>y��HRc)ȓD�* �$?Oz��L�r�:M�\�H�| ���� d.���'�.���Ǒ����r�Hp*QGz�~RQ$X�E L���   �  �  m  �  a+  D7  �B  iN  X  !_  k  �s  6z  }�  ׆  �  a�  ͙  "�  ��  ڬ  �  \�  ��  ��  '�  j�  ��  ��  6�  ��  D�  0  s  ' � �$ + �0  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c�>���I ]JP�D�B3g�THD��J���&"Q�"}b���[�9g,7aj,˗��e�<���C6p��-Ҁ��#��k��a�IZ�tR`˘/����6Rr�����1$�T2�jǃ%��|	���2B"��P���0<��4�O ��Q���u�XqR��k�<���"O:(Q��W|�%�_�(�xS�D��,oR�)��<����䥹��j�i���O��hO1���D�ԯ(� ݐUH�$w��pa�;|O���ᦁ<V@)����]�#S�d�.��'Ҕ��cg�O<6���hď�A(��a�8D��:��7CΰbÌ^���&
�2:*�?��d�	-��P��HZ�S�-2V�a{2�d�3Ђ��E /�<m3խ.W������Fx��)@�A?��c%	�,C�R��R�A,S�!�d-x<=Z��� �T��#�x�D5}��'2�ICF�_V��|�t%�8�X<�
�'���g��8�D��An�-�� ��:�x�$s`h{��F
��!b��1��O4����ю L�ZP���D�>�dW�N$!��f�T��J����a��DqO�=%?ysF�o�eGd�>]�$l��',D��;E�p%t h��3L���Ff-�d8�O,:��E 9b�La���8r��E�OX�L5a�T�d��*��٠�N�-e!��W	$A���-{�X��v���]1O�����8z�ѡ�R;#z1:�(Y�]!�Ċ�\��$�#i����]�^W!�d��!����"�HPm�u ���A!�$͢Qa�����irm�PNJ"uI!�Ք\$����HR�e�$�Ԣa{bKʦl>�Jd�2@b� *�p��"�S�D���J���3m�}���;p�)m�耄ȓE��A�;q*J���ߢN��p��	;q�O�͒Ю�/c�21'��Cr �p�"O��kR-{!�X4��1j֌3��|�)����\+�DQ?=���J�G�QJ~C�	)>���; K�S�80��ر+�^�� �DL5�Pݨ�@Lr,�9ЍL9	7!�deJ]��E���:G_�#Q��G{*���{B�
�4�� �--l��[�"O�T	�O�r�����,?V)"O��(�M��4<����E2/�2�R�"O�	�q'�4ȼ� �x�����"O -�U �o��(p��:.-xԠ"O\ဦeG�TZ<�'�aS�"OT���a��e	*�v.|��iC"O����PѪ���lВG0��:�"O�I�i���6a!.�?Y!@����'Wb�'G�
G,�0�������0�'�jS�o��;MB�hc�ڡ�@�Z�'�f��6&eR�,cFǶL�R ���x�آ=��e	����CY�rᆜY�*�V��m�ȓ�
�8yZ��vEN;�Z%y!�)���YfF��)]L,(��EP�I���&D�����^��RRg 9 �0�Pr,�>���u��P��<y��hpÊ׿Ian��ȓ-����c��`�(c!	�D=� ��S�? ���E��65�^�:��������ȟ��C�,��$ڪ9 b`�3^�e�B�',N-o��$D���$D�
�����.Ew��Q�Ðg�B�F{���'�X���C�4i�Y;Â�'1���',���0�Ȅ
b�z������K>IJ<����� 3G�ϻo����cڢ!~v��"Od��2Ӑ6��tq���Lt0��2"OV��t�܊���Y���+Q�|B�'V��t�'qP���l��,�(LA!��U*M�w"Or]2�m�X�,�H�$������>�y��9ON��T�̈x
,��҂�c���9�"O���+�`m܉�7$�F��!�"�i����=Y��S,;�Xr2�!�ju�t�Sc8��%��RtIyYԭ����)qH$d�I5D�<�bN�I?�E;@�Ϣ[���RQ�3�d�O�i�<����Z��T���J�]	e����4�C�	�7�AA�@�/H�!:����9�?9N�[���$�(� �I}�ԅ�t+Q��!��F� �����G�!?��1pQE\=Y��ĉF؟���
D�~3�����s�b���x�?������XQ�:I�(1�PM

C�p����82C�	2[z樲�Kز'�h�h�Z�3\��I��!{B��"�9P����gĹ'Eڠ �;E.����qx6��3�O�5��tsaзeԁ��5Z=J�HNN4�P7Ҷ�����k?��	9{��0!�A!&�x�Ny2�'Ʋ�k��-8�`ܠ7 H6|0��h�1O��5aߢV��a0�F�u��!jw"O�"���%*��u޲R�
�0"OrL���OǪ`�.L�u��h�"O����B��v� b#%���B�i�ў"~nZ��Z�윉	�L��B#�elHC��,g:���o����ۺ8C䉔w�	X��Ĕ��]�E� ��B��7~5�7D_yْ�j���B�
i�ԁP5`ڽ?x^�KT�Z!�B䉸i
�:A��X�*��A��|��B�I�g�Hi@��L�0�lH�,O�T�B�I��Uc���q����B�HtB䉞$PL�A�Dɕ'��	�!�SB�	�y�d��B@"_lM����3(
B�	�3���A�d�7G�0i2��D�|�C�I�aɪ��F�_=[�*sL�c�C�I�f�����,����	j��B�ɒ/~�p���q��`��&ٚB�I�Ba�1�>BP̌����G7PB�I5%�ph��9�la�ǯ��m��C�I�O& �#V�ɐ�~��̏�8�B�I�@����U(~D�ba��3:ˀB�I�Y^�j4D�/&�>�2I��.�dB�IW[�݀ Î4����ɕ�q�BB��3	.Ȍ���W�4��DY�H��T�LB䉨R��L����RãФ"+ �f"O���l.kO�%*��_�:�x!��"O��0�D�5X�1ybG�a��X��"O�����U80c3�s���PT"Oh�̊��>���a ~�8�j�"OR�YK0���:� �m1�D"C"O2d��ِ
�"�B�/�	-�9�'"O&M00��p>�b 	.S��Y*3"Or:�K@�=������4_
���"O褫%KC�UY�o������"O.���MJ�(�J Ǎ�p� �1"O"�#A�Șx����P�GHK��y
� FP�%J�,�8! l37H���"O�[�P��έH�+�0v8�"O�m�C?t�����3`,B�"OVWɦP,�4�&���P��x�<v'��C��T)��ћx戝S�kL��D�Iן��I��h�	՟ �	ܟp�	� z�*I�#�����W!�=x��������$�	؟������I����ϟ|�%��"��e�#�]Gr��^�����OR���OT���O<���O��OV��eHb91��M9z�QFŏ�.T���On���O��D�OX��O����O��D��B�ޕ� 	.?�(ũa�΋b<����O����O��$�O��D�O����O��Q�C�rE���b���gFQ�?���d�Or���O�D�O<�d�O���Ob�Ĝ�Qs�4y��F ����j��JL
�$�O|���O���O����O�D�O��D �
�2��/�8Ht�=[���?[qh���O���O����O����O|�$�O���E?x�&��Ê�XDB!fM�YCJ�D�Oz�$�O��D�OH���O��d�O����~���	�zI�R�%U�a\��$�O����OX���O��D�O6�d�O����@�X��G��}�Ɯb���\���d�Od��O��$�O,�$�O����O����bk�$��ȸHW�$ �����d�O���O��D�O��D�O����O������A�
r�8���x�R���O����O����O����OF�oΟ��	�6�����Ѱ��j���L�*�a+Op���<�|�'(l7�%K��|сn�q�@�k;}OJP�q��,#�4�����'e��Fm��
w'�&7���H�lX%+�B�'��SR�i�	�|R��O*�'$���#"f�u��_�P����<���$,ڧ5�j��0��|ݐ���{&��ra�i"�)�y���Y¦��t"�P&K�Bڎ]�f��jX���ڟ������h�#�M��'�D��ǈ�S�v�Eo�Ev~Mk�'|�D��Xt�i>��	,5`1*����Xy��jΫ��Icy�|�Lq�8pb�dJV:�Ԇ�$��<#�咵`ܤ⟼ʯO����O���~}R�\���2fX8SU��������O�$ѳ�<1�1�� ���1�h�D@:4]A�C�J�8p��Kw�ʓ���O?�	�R�ni5.U$�֬ȥ+XUP� �M˃�DX~BDq���SK��h����:Us�P{֪G#36�֟��I�<�R��Ҧi�'���?�2�ȚQ;�W�����H�R�'��i>��	ݟ��Iן<���#���:W,הiV��P/p9>d�'�7� !�r���Of�d+���O>E��l���5���L����@e�o}�Epӈ�o����|����:��ַ?��̺��
58Xd� �P�4p�B�̊�?�P���F@���u��&�ny��Ӫ7�舥(Aq|Q`�7/e��'���'�O��I�Mk!��?y��A���,l�MHAe��0���������h}��j�n��MSaI�e���Η�Lc�1�
4p���4�y"�'��F��?�1�P�l����y�V�. �&5��B��<h���B�w���	�� �����	����j�Ճ4�>�B���ܕ�B�Z��?A��?Ab�im(	��Ob�guӒ�O,�+�7�xQ���p�����Q�I�M�5���4+�?��֙�H � V@F(]
�D!$
�馉�0d�fH�'�L8'�\�'��'���'���	գG��|���J� ��Q�'��Y��ݴRuFY3���?����,z�Q�f٫1��)�Ņ�TH���O��'�R�'�ɧ�t�'��� g��("�ᄥF.�.p*��p}T�������?�A��'ed%�hJW�I�&L(S�&B>�D�P�`�I����	ߟb>ɖ'ߌ7-=`�QD'���"fb GUbPA�<c�i�O���'q6�xʁxa�؜����<�$m�9�M[e,ɳ�M��Orj������<���E�S���[�m�>j
��c-B�<1-O����O����O<���O�ʧq}��x���!Z��uQ�*R�B���0%�ic6�id�'���'���yҫr���q�^���:�^��0O��I-.%lڃ�M���x�O����O+�id�i��d��{IE0F�ɝn��Y����2'�$QU����*��O������5����P������5�O�*ax�KrӮ���<��l�r�A���4��h>3L�����e�>�f�i�7��c�6r(LcPG�!O@f\��L�7 ����P�m�i�� �dy�Oˠu�Ʌ>��ݝY%&+#����D��ñ5�'���'���s�ոDM��Rlf� � X����V"ϟ�S�4{�`-,O�n�z�Ӽ�F]<L,H�6�0����L?y���M맻i�,�!�ii��>]n�$�5�O��}��ڬ=��x g�#KӖ���,U�cyR�'���'���'�gli�7��ѠXyvbJ�ؘP+O��o�*�.��I۟���F�s���a�_B�!�a�#M��Hk������ͦ��ܴh���S,U����+�\V�褦�7k�t�  *����'ج5�E+�����"�'#�my��ѷ6����Ν�A�M����$,B�'�r�'�b�9��'�剼�M���ݔ�?q�l� 5<F�0��]�
�cPK���?��irS������릱��4SΛv�G�D3�jY��z@��>8`P��a���	�4�'"GC���xy��O� �܂nA�+��qh��I�HC\�{��O���8���D�O��$�OH�D�O���,�O��  h
+�t����O�v��bT?O����O`m��C���IƟT��ϟl����`hѤ���8!S�I�C
�3���?�v����4q�f�O��"e�i��h�>0iQ�D�U�$a�ȭ��x&�� |�{��'���'���'��OL(95MVR<�Mc�'U?]"���&ብ�M�� 6���O�˧U�ܭ`W�����ҁ{����'���?Y���S�F�w� ��X�p'�p
D5E�`ygLɘa2����V���5$d�/�I�Tg$a�s۞��֣Ȕz��B���M{�b֏A�1�Չ�$H�]8��޴)(�8,OJ�l`��N��ןLs��� ٬�U��(ȒA��\��. �|�o�<��O����%�O�(�'��m 1,��<��Y�"K4`�ҙ'��Iȟ��������D� ��e��A�S�{3B�JG�AD�7-�v~��D�OP�� �'�M�;S�,�-u���aiC�>Ȍ�0!�i�7M�D�)�S�Y��l��<�P^�>A���@�ֿd�Lx�t�[�<��Kpt�䇧����D�O���Z�r��H�$��%O*�Zb�]>����O���O�ʓ<����҂N�'�2!��
��@�@Zn�+ i߇a�'Q���<I��M�R�x�	Qs"n�רX39�Ti&��"��$Q�+���O^�G���&���E8�Ց�	��ː1�x@�b�O-'���d�O���OX�d>ڧ�?A�e��6L����A�w*�s�)�7�?��i���1��'o�nӌ�来J� l"�nY�Z!��J �Dx��>�Mѱi �7� 7x61?9@M� �2��
�Z钷��T��q�dW��e�J>�-O����O�D�O��O���F� sz8X�� N�=a�ă�<ɒ�i�*�S��'���'��y�햾q�=��Gz1�#�O��
�0�|���i���%�b>A�fR.�&U����:O��Ab��6?�)nڂ�������~B�|�\�`�S�[2��5H8_Y�]q�E\��4�I�����ݟ��[yB.r�$9ؗ��O*{��V�X�h!#W,@��#���O�l�i��
�IƟ��i�Er���p1����2N���c6��a0mZy~�Y���-�ӎ>��O���#�ZpV�.�6�q�&б�y2�']2�'22�'�����>s���P�+4Y����7&�$�O��d[ަ�Cb�b>m�I��M�N>��C1N�-�%IĜ\�.I��
�im�'y�7-Iڦ�	K��l�z~R���4M֠��_-88|���˄@P��WE{?�K>�*O�� �0�A#zhT�fE��cb�9Xc���(��	��ȗO����d �dp��%D
t�x�c�O���'d|7���L<�O�NH"s`S�����T��&T��	�섿2��$�s��i>]���'=�&��j�%QF���	�"�r�Q���$�	�����ȟb>��'��7�""�,U�ƤW4|b"<$$ڬ&� �G��<�i��O0<�'�7mˆ��V�șcR.m�#X�6ilZ�M둎�MK�O��bE)����c�<�� �<Z�&����ƒk<�x@�<�-O����Op���O����OL�'?V�2���-c�n��d\n�.���iV���%�'VR�'�O\R�t��l�T)�q��)�p؛d�P�Z�P��	⦱;J>%?u�pj�ɦQ͓����nlMXpi�+	ol|̓}�\ fA��l%��'Zr�'�XɷL�!_�h��S�|tn����'���'��U�Xkݴo�\��?��(ⴴ�򫏢w������0H=6ոJ>���\�ɵ�M{S�iS�OT���A=a�t#�g3����b��(�BϒtC��Cg�X�StE2��ʟ��u�BN�����Sv0�ECٟ$��ϟ`�I��\D��w�b�8w��6�|eh5��'7�x  ��'ô6��/F���D�O�yl�p�I��^, �`b��X
	Js�+��物�M���i��6-�4��7!?!��"]Tl�)$0s�%��̊�Jb�!� 	1�X�YI>1��?Q���?����?	��?�3 �NPV��@�"P�::U� �?	��3P�ܑM�#�?����?I��i���'"C��hD�J��ɷ3������_�ztq��'H�6m����c/��?��O����q��ͨ��h����Bk��2��*"_��HV��<a�/��n���Z	����dRD�ɐ�Ĳ
s�#�DơR��d�O��O,�4��˓N͛��ď|�".S.9�1�J[�6-�Y� ]6d���y�B�� �OZo��M[��i�H|9��ثoЈ�;B��!<�y��`��<w�v�����7W��d���߉��)��J-8���48CPĢb�q�|�	���I������J�bZ! ���j�oz����#�?���?�T�i�p�+�OA�p�4�O��B�S�@��'^[�x"čJq�ԟnz>�!cLZ禅�'[��i���&<��(����hެ��s,Ss%L�I1x��'#��,�I����ɚp^J�{RH��D��0 D �5���H�'56-b�p���Ot��|JD���cR&�6O�+h����"-�t~���>��i)�7�YT�)�rDƫ5yTT�Q��z*9;��--G���'�����-O�	�)�?1"�>�	�za�Y� �]B�~�K`��8�:�$�Ov���O���<ip�i��T�AB�\�4�G�A�[����"�ܳ'��'�F6M2��'��D������65|�	倝�r�P5���ʜ�M���iu�a�ֱi0�	�4��)e�O�P5��� ,5 �O#\�0�J�����P��p<O���?�4A��?����?���?�'Jg��	�\��^�7$�$,8����i'ܝ��N�=�"�'��d�[�b�'�w�%�G���V��d��iA
q�X(ڰ��(�m�-���қ�O��$�O��u"5�i���Ӭgo�Hp  �?G� ���O̻6�d����f�F�O���?��T�D�x��J�nE���;@�������?���?�,OԸm�{���	���	v��m��.��2
p�w"Z�,��9�?)`W�l��4]d��K<�$Z
��-{ N�����ՋPx��-.�MADAԈ��m&?=I$�'��M�����j���-? �*Z���覍�O<�D�O6��O쒟�蒠��O��d�J��p�ˊjX����$�N���ЦyS�j�П�����M�����$�O�پN��;F�	�jB��c_�����ܴj���Ub��61O����1G�ё�'B��x	�E��T�Pݑ���	/�B��m!��<Q��1Q���V+�d3F�&�J�T�	��M���L����O��?���$�tH��
ڒ=06��?��D�OT��!��ɑ�#KN���g�~�:�1� I2^����i�v˓%ɀx�"��O���O>�*Otd����bH^5�� 3HQ�(J���O,�D�O����O�ɡ<�0�iZ�2��'j\Is��H� p������U����'��6�.�����ݦUX�44���m�L96��4o"� ��FM9��Ѫe�i�I5���՟v�������YR�x�K����@��˻l�d�O��$�O����O��$?��D]�b�M�n���B�ܠ8s8�	��Ɂ�M�g ������$� �cN�a>�Q 	ץtr�X�@ݒ�ē[뛖!m���IE�7$?yrGф%�
����Ѓ=�vdZB�(e�`��bh�O =�I>�*Ob�$�O����O^�yv�ʿ!�:PBӨ��Qu��C ��O���<Q�iRΠa'�'��'���+D�Y��iX�~4)K@��V���N���퟼�	u�)b����g\,
f��=4�ʰ��w*<�zWI��K溼)O��ߥ�?��&-��Pb�2�O�my�S����l�!�D�ڦ)�@��'y8i�/��1*k���	�'L�6�0�	��D�Ʀ���䔙.l�I��"�y�X�V�O�M#�i�>���i4�	�/��1��O�Xݕ'�#ъ2'#� *�Q7����'����,�	�@��͟|��H����zҔ|K�	Qüx���'*ڤ7͌�w�d��O��3�9O�ozީ�QO9��1
��F�֍�f#���?�۴>�ɧ*�'�"��X��M˞'�`�eF�=x�cu �!�MÙ'a��h!���R��|2R�|�I���ZB���|��A��#�w>����l��\������	Zy"�z�v�j�h�O����O�P��N�6�ޝ��M�w��	)�//�ɱ����=2���'���)V���v
D�p7�שDf����O�J��6t�^ AQ�;�	�6�?iQ��OH1j�	DLe�!�-��� �I�Oh���O:���O`�}��w^q���(r��$;6�eƌ-b��=N�F��a��I�M��w�jQ0H�pW��i�Iͅvs��r�'c�6�VئuB۴"n����4��D�=�ڈ���h 6E�pET��n�H
X����:���<���?����?I���?!Wa׋:���������a=�����=�m�<�	ޟD&?�I�B�uk!��(9���{�%C8�!P�O���OƒO1��h�`-h`��/-�`W@
� �H�PV��<��V#�����%W�!�Z13�lşZo��iꍨ!FJE�%��F�Ҽ2 �O5;n�&�O;L��1�T��.��$��b�+\�&b���r�h���D�mĸ;�E�k�xxp�Bj���[<��A��l��r��y�� <������ôp+��#vϜ�UZ�a#�Z(
��%I��B�el+����Q>�5���T3���7"���E�5%���9�(D(	|��"�$W�!D�-���B��ț�� ,��d:��z��K%j���}"�
M�I�z��B�� lжH�3�ҹ�&�sw)�O<���Ic%����/Z`���O�(ݦuo�0�I̟h%�4�	�<9eu?Ƀ��6|����b��`u�]}��'���'^�ɀB��m�OZ@*0`ds�Y�G�lu�'-H
��6M�O��O��d�O��S��8a��
�JU�~Y������
]�6��Ol��<Q�E�3��ן0���?��׊��`���^ ��W��60��x"�'"�%͒[��|Rҟp��J�6G���y ��/Ǽ���i`��,	�j�#޴�?!���?��'��i���J� &��e�������B������(#7�O���O��P��G>d�4W�Vz\�޴Z����?���?I�'���O,�.����o
?_��2���=s���l? �4A�?E���'�^�«�5d� �
&b�(��@7Oo�H���OF���r�v��'��I�`��,��9�����I�Ч�G_��>iwm�Y��?���?��Z� ��z`.ωLEz	��M"aj��'��bŨ>9.O�D.��ƺI`ԅ�^�q�AM3H��q��R��A��(�	�T�I�D�' �< ���r�T���$ܧ	��sPKױ'!�����O�O����Ob���I�\��)Pb�i�J��Z���<	���?����W�R�t�Χx3T����o���\9�P}!պi���П�&�p��П
"�Oi?���*GF�dba�Jm�$ ���d�On�D�O.ʓW@(�&����T���ޚ|��E$� Mv�m�ʟP'����ʟ��TK�|ܓ���S�O�-��Y����8`��m�ϟ��	ry"�<`	�����?�� ��x%̅.!���I�
s�����x��'��Mπ��O��P $蚰�πB�:�Ju
ټ6&�6-�<������?i���?����.OkL܎�j��@��
=��bE��#	-��'⠝K��O��Rh�!n��0l�b'��Vp" �i���p�'��'b�OT�˟��q1%�V%^��-�W��,V�)0ݴ) b�����i�O�H�b�'c���TD[=k1(A��i�����l�	$J�&m#L<�'�?��'�v���dX.���8B#$5��{�4�?�-O�U31$�[��'6�'���3��δa'���wٍf��7��O��r���P�i>��	s�	�C�,���I�m�����b0hO<�����$�O�$�O$ʓ':����-0�t���&RE�yb�枂Z�'���'��'��iݽ�Q��b@`�ę�e(Q��k���$�<��?�����$(yͧe�X��@�Èy ؼ�Vb�6�F��'��'��'�I���=��!W����Ѕ\)��q�e$�;��,�H<�����d�OZ�����|���W�I�l3�2e�'+��::�`�$�i��O.�$�O(��S�A[Չ'�88��#٥l��W��/}0��ڴ�?����$Ϥ�I&>��I�?��R��l��\�'���{���_W�6͵<����?93넶�?�*�����k���*l.��U�E",�4\��iܞ	��	�p�t��럌��ӟ��	�?���u7Qp��+uC��p����jR��M���?Q����j¨��<�~*�k(TiG�A:C>�f�RĦ���kDן��I�|���?q���I�I���So� 9��� E-yx��o�g%�Q�׈/�)§�?)򫁌A1P�S�Ĉsk\��%�g�6�'x2�'�>ћwB>�4�r���O�Ũ���)Vd���\�$�7�Ҧ��������@�B���'�?)�'��ev�0��$\04J�U��4�?�Ugݜ���Ag���Đ�J����c �f��CW�U�H����'��d�b���d�O<�$�OZ��h�+4t�e!EN�}j�iQ ž6Љ'<��'o�^���I۟�A���'L4���4��U����%�*y���Iwyr�'��_���� ������-x7jIߐ@2S�I9%��mZ���IB��?A�,2I`5�צ����-@uxuA��Z=��볅�>���?I���$@���$>a���K�}b0	��F=W*�s�M �Mc��?A*O ���O04���O�˧'�L���,D3��A1��
JB�h4�i��]�T�I~��	�O2��'��\c��ƛ0�vq	#ރs�l�CK<����d˙���}#�l�&B�,P���##��)],�l�UyR�G�TZH7�YK���'��$�4?Y��G�������jZd�!��]æ�'���'���'�~��B&9U�t��ё�f���jѝ�M�� �?���?����j)O�&9
%��P1K��p�w��K�U�ܴff}ґ�d�S�O,I�-[��d��)w֩�^�/?66m�O����OZ5�C�F}�T�0�	u?�`H�	F,(+�
������A����%�DC@b���?A���?s�Nl	T9Zd�}���r#�	�U���''�9#�>�)O��$�<���ӶEǢZ�0�2��R3�x{vIզ�	�R���� ����X�����'���J $�e-8=�5��%(���"��I��듅�$�OV��?���?���z�J�N��}˴�-~k�H͓��d�O���O����O\@�Ӌڦ�Dn��I��P��ūnԈ1`ř(�M���?q��?������O�왗>�k�T�.��$�Ԫ�q��)�L�*Q���'���'�BU�̠�f߂����Oklȋ]���8�i-u줉 �.jf���'��	��T�����S��d�X��M3 �3"�Riw��o�R}�`��6��Oh��<�r�Y
J��矠���?�a�� �%��h$䒢p��Ң������O�d�O�-"�4O~�$�<��O�0IS�P @�� L[�}T�ڴ�����l���	����S�������E��.�|��
�(e�]%�i���' (���'����<�����&�j�
%�P�HXޘ���;�Mss����v�'.��'���/�>1)OFq���-�����h:&+���q&`z�x$������i����n8&q�bG٩�t�R��i�R�'Vr+��Q�������O��	w+��P���R���q��7-%���'�?��Iӟ`���o"ܥ;�.W��xy����O��%�4�?IU��S�I`y��'��	���أy�B��7cD ���d/�d� �L�4�̓�?����?����9O�hY�ᛍ&�F�) �~�
�av�Ū1N��'0�	ӟД'1B�'M�n2f��P�G�ڣYt$B�I�5%J�1�'r"�'���'�2W�@��!������� . �X$	)�b��C��MS,O����<Y���?!��
���'�P�6e���NE�0�7<����4�?y���?9���D�4��h�OvR�T �tN)g,�1N�h7-�O���?q��?a"�T[�z����֍Y
 ���Nƍ,���mZ��`��{yR!XQ��'�?����z�M�=�*x��T�8��ǡS�p�I���I�����L`����yBџX��n��Mm|�c�N%=����C�i>�I�I
>�Rݴ�?���?���'��i��@.ٲ[�b���ʝnV�(� i�����O�>O�OZ�>�P%�Ϳhc�嫣]�n�&�hӎ]�����1�������?])�ON�l� �E�r�M�k�Z��@n��8��a�i����'�'_���ȉn;3F��+\�S�-�H��en�ğ��	ӟ��% ��D�<!���~�K�693�%^�d����Ms����d_&/s�?������	�6�H8S�@�0k��ŎbIB��֦=�I��dѭO���?Q*O����X���l�8��8CF��9�0�H1[���S�x���	ʟ��	����I\yR����ll�*<5Nz%�tF��*	���>1*Of�D�<9��?���a�������)i�2���fu@���<���?!��?����DE�=Vԝ̧fT�<�JՉ(�j��H7i���o�Ty��'U�ԟ���˟���s�\y4#K�_��B����d
��s&D�M���?)���?�(O�L�VK�r�T�5���VO�e��f��2Uĭ u.N���_ǟ(�'*��'�bB��I��0��&=�>�t�)pj���&sӤ�$�O��M��!�Y?��Iܟ��L
�\�)gbr�R"b]�P����O���OP�E.W�)���?1�uH���ճQ�H�p�:�b�/p�L�~�8���i��'�?��'q�� x_�`2M�&�lXѯ��H�6��O��D��zM���8��=� 7ur�;�o���,
���X�$6�_46̬@m��������@�����'qr0`@��V8���$V��� �%a�J�1E�O
�O�?y��ulN��o'�E�ǐ�g�֐��4�?���?u�.��'P2�'L��V�8r�5S�a۫!�f`pc(QڛV�|�H��������V�'p�̓VA.3���,�0g���Cd�,���+~�`(&�P��$�֘F��ae�*1&��ұ�e�l�#�F̓��d�O*��O��e�Q����0!*�X�O�':$�jf@�%Y�OX�d+���OZ�DL&�<�*tO�jԢ� C�H�v��q;O�ʓ�?�����'M�<�V2�����ʗ���!J@I�=����Q���	ڟ�$���Iڟ��c�q�tauʀ��j��OS�Bf�)@��5��d�O����O�˓��D�f��d���7�l����3�u(3#	�t��7-�O�O���O2����<�0�B���#�8�ad��@�7M�O���<ђ�՚*"�OGb�O�B ���O��x����P(f$San�>I��?I�z���Exrޟ�-�JƏnZFd��_�a��i\�	�\��ش\��ȟ���!��dT6,���cQ6A\r�I�r}���'-l�%6A"�|���ON�=���iwKW�S�m{%FR7�M;b(P�'���';���=��O��Fꅸy ���W�`�b���æI���ß�$�"|J���hP�A��, ���^
�� b�ib�'�bQ���OB�$�OX�I5j<Mx桅�z@��A�B=^Z�6� �䗓m��`%>���� �	O�ݰ��A��<#�I]�4 ��4�?᤯ǚG�����I�k-�шg�V�'t�� 	?���`�����d�O����O�ʓP���c��B�N!g	�d4� �f�<rj�'�R�	�����I�jxhDy%�@�x�WD b� �I�����(��ן �'��X��f>��%k_99	��y ��(n��)�CJe�r˓�?�/Op��O���T���׾^2��YB�_H��L�,���n�ݟ��ɟt�I|yB���!����?�SG�?f� `�ƛ�^��i�$�L����'/�	۟`�	�T�n}���Oц)Ac�D&P���p��սQ'<qQЇu�v�d�O��D���tR?���ɟ���\��U-[qQ��T��2��h�OX�D�Ob�DM�r�$%��?�Cg�]+:�4h�6g۔e1�J��x���C�6�$�i���'���On��Ӻ��b��ցZ%ʞ�|? )���������D�&	'��Oz�-�&/J5��8U�ݴrZ2��ѵi�r�'��Oż����8<s� �B�[�r�6eY�-��Anږ9v�I�l�'j�b�$ h����k����\�U��.of�m�ߟ��	ןL�P�̲��d�<���~��LW���Z�
 $#lڅ#�Ɔ��M����?q��W���S���'�r�'\=1��!7����	�R�n����d�6�d�2:��,�'����ĕ'�Zc~��"�&wХ��3`H9k�O$�3�=O�˓�?Y�����O41S�J���p�������2�'�J� �$�On��ͦ��	`�I�����m�)�Q�)����qk<e����lW�bz���?1��?9-Oh��w�R�|"`m��{���W>~(�e�}b�'�|r�'��;����� `�0�J�+�:�Ñ`N& ��ȟ8��ğ�'Z,9s�K?� s-�A[4d԰(]��q-��ll��&���I���$�IHvƔ��#0+2� ��0A*��`G ����O�UA��+wA�ܸ�i��`&?�̻}�0G
O�F���
´{$a�ȓZ�zLbP�Ï>�xz��߹2�.��EG��*԰�a$p)�ճsn�Q�H$��)@11��b�[0!�~<��
B/1� 
A�YAeG��:Q�Mp`��*m���ӂ�nLi�Pd��F�K�G�3�\��)jʑ��j��L���!tET�z�(40Vi]�aD�`7��p#�a&��P�,=�� ː	��5���?����?y7��d��';u�0y���C�l(m8$�Ǐ7�	Z�^>I�r���t2�b>K���`��� )��k��V��sG�U!<vD�

И'Ǜ��
�B�T42���t'g�7=�x��E�'T�|�F�_�d��q���O��[�&��i>�E{Z@�K��/|ɞ`:��T�BQ^(P��� ���D��jQH���\]��$�Õ�l[���?�'��Ҵ��"dkt٣Ӥ��.s,�!�?J�
���'c2�'���uݩ��ܟL�'L�������/n�*�� "ר��$E50T��@O�5L��	� بh�bG��\㠅�20�z؃f*�F�A�(�-9;��:ϓE�}[ A+u.�ؚ`dK��T سo��|��`�'��OD�գN6$���Q�恜l�#�"Od,�`^�b�t�`C��R�ZD��~}�R���　���D�O��S�%�;�^  �r�z4:$C�O�d�`����O$�ӗ��q�c�b���[���妉(��� )H��U��G�j�Ad'%O��fMښoP���!� LD6�#]`��'�0I�D+�"�xb� �?����򤛉b[����G�1�T��@�1OR����v�̤�G��T�� ;�<5!�dN�E��fJ6V��r�	*���9�m�$�'g�͘@�>���i�/b���8�N��%�!|���e%� W����O"X[��G�ov>�q�dS��R���|�/�:���/O�l�܄�G͎�*�D���>��	ԇ ;�5�I�'u*]p��0Z�J`P�O{d�3�l�<s&��Ȑ�IʟD�t�'͐�$@��	-��b��t���'��y�jX�| C�f�kK*�pÓ+<���A ��!U\�(�dE���Y�v����M3��?Q�|�l����?Y���?1�Ӽ+  ^�����uV}��R�5�xOr�u�E1g1��'��1j�mR�;80��Ɗ�l�j���z≆,��Uz���|�Q�3P�e0����l���Y*�X�7�����I pVu�)�<Y��l8�={�NC^��Q�Pi]������'G�EZW��'�!��B�Q�TP`�O��EzB�u?.Oh0;�F٭7����*������k-\2[	�O��$�O�������?I�O�͡�*�Wp�*A��`h6A�N��O�z�bG��s8�`j�- �BZ�-�f"��\�Q��h�!
��$��ӹWD�|� �=t,9�E�%ڰ�$A��F�q���?Q��?�)O���7��3l�<C6��'bJa
a�HdBB�ɡJ�R����%b2U�4�?�Bc��9�OʓQ�kc�i�B�'���pG_E�A�RH�,M~��1�'a��/��'��)�k������F���DW$=��es!��?J���cĘ�g0�x��ˆj����eI~rh�"Y���{�%XLZmk�I���p<���Ɵ��Iߟ�	���ـ� �v�.�dDT!� X�'{"��S�p�z� ,�8s  ��-�7"�>B��:�M�Ga[6X�B�hD��#0$��ʹ�ؔ'#8�s&Iu���D�O��'����`���!Mp�dah��ީ;��R���?�w���?��y*��	�I�ȸ��j0�|��R"F��''��ٍ��IفL��UDր�	��Y&`k�(��Iz�S��q�zԠΊ7��ٛEɥQ6��FҚ����\W�twk�#&e�h�ቘ�HO�UHC���Q_6��B��f\ے	Ŧ������		n)��i�ϟD�	����i��t(��W͚�I,�?8N�3���n�W�=�牷o/��*�˿a���!��+
�����9<O�j���	,�dd�+���d���3�ɼ�����|2jN�/��C�&MUȍ�5�� �yb�ݧY�ꔬV�@�H���.����ĆR�����0n��r�1R�f�!AXb�{�iA�p	U�Oh���O6���ͺ����?9�Ob�$��JةN���"̀jN�hK�e�=�L�&J��*�Ԝѕ�'���#���"}�,\�7����<<Sv�gjԩʵkL-zB@�9��'k֩�@�Y�`A~�!�TF�!O]��?���?Y�����Oj�4h�Z'�E;B�'�T���'D�tYeL<~�X�R��,�P��5D'�ɡ��d�<�q�ԟi&���'����Qȍ�Q/M��0ؑ�����'I�5���'��'Pn	���R���X�FMP��*�s�������61g8Ѻa#�)i����%ǀ8�T�FyrnH�G�U�B���Y��qK"�,�b��_ " � ��0�M^$E$%DyBdR��?A�I֛&�'uƽa�	�2,ʈ����1<RyX�W���I͟H�	]�O�`���F�_� �)#����
��x��yӖ�zdLN�|@d�D�J�T���	$���I��E{�-�e$�Ĉ	�*�W`�	�y� �A�	Q4cR4MD�D���yR+�D�6ًC���I<n��%4�y2F�-�h�3"��=`R�,�yFƝq�$�q-�.�h�����y
�  I�TI�6Q�D�/*�9 �"O�qy��X+$9��-W�����U"O��˦�TO��7��K���g"O6�1&��5]oذ��a�$D�A+�"OJ"R�ȷ%�J�i���4��Q�"Od��HPM��p�5�C�T�
�(�"O�,R͓�L{��*iM�QϜq;t"OA�g*ӄ$�pb��5���&"O� �ҬN D�R`1h6c�4�+"Oq���6�P`ӁΉ?r�q�"On������7W��ak�(%Xy�6"O�1�e�1����A6�&y��"O�h(��C6V���A�iQ�7��� c"O Ӈ,Z!A-��q�Y�e͒��"O
9#,�?2,MZ����3!2���"O m+R
	=I�ӥՁV�z�"O�����څVN��aQ.	G�j�H3"O� �禟 Fx4����n��˶"OR�У��wf}��� Bd�t��"O�T����$��8@��5'6��7"O�Z�T4&������X�$T���"O��2 ��[���qQ�W3xlBY!s"O�q�kC(0D�k2�D8I LX�"O�\�MO,"��HT��%!�J"O$��׆D��|X��F �fUh�"O�uy&�?ZՖbDF�Z�Pi�!"O���s�?WD�-�ज�H�A�"OJ��6�����+U��{$�e�"O�$:��� hʈ8�CыN8�"Oi��L��(�֬��j�Qh�"OZ�c�1o�  � ��^��T�B"O&�Va�|�`��q
���Zع$"Ol*F`J�Q���&*T6TX�@ "O���mk���TCX��4"O�h  �4^�0j!O�3,)�w"O��@�*+Nl�Q���F���"O`a��܁n8
T�@�< P=�P"OV%3f��jE��!�1����"OR�����=��4��e R��,�B"On��")Y?/L��bEeۊ!��U�P"OTm�V�_.>��`(�ĈK��pcf"O9����4o=�Q�V"���""O������Ŗ�%#L)z�l �%"OFdQe���(;ri��>Y6���"O��.��y�~�`��f������9D���둅�LY�$��kmf�Sd:D�0i��^�h���1&*�+��$��7D�T� ��<Qj�q��4�`\�7o7D���^�t#�m �#��foJ�j@�2�$��&�J���^�0!#V���n�<Arg掍�a� p5�L���љ8j�P�W�o���iǀ�vh<�3��I[��""�+G�<`���T�'��i���N2��O��8�QJ��O(.�{��M.^�"U�	�'�0Pr5 t��0�A� [�$ �O����䑛J�1O�>��*�	
�F%� �7"��&�<�H�����(����@�{�֜�'�,�u8�xbGUp��P��	Z}<A��&]/$A������#MܼO���Ǖ��O�xAF���tܸlB#��TLy0'�6�2uKۓb��� ֎D�.�p����,���k�J�%���qB�y��Or�ҰNN�S��yh��YH�'0&cW�Һ|�,���ӈN^��>�0���W6��@�M�
k��?M3Ɂ�: ��q��Vp2���3Q�9�h�	P'HH�0��>���}9���]�(Z"aҍ	���c̷C\N��рR��~��4�g}2�O+TR�y���0۪-q4�N��Mk�R\�u�nK�e����wJ��#�LIhEpe��|���FY�rqz�a�!�H.Lt�=ɔ�^w�:qˑ�� R9Q�,"v�S	EXa'Ő�6-�A������ɣs�\$ji��T�ks�Q7 ďq0�Aq��<~QPa�5/�z~��!<"�� gfݩ�טO̡z�D�,�����aQ�.��]�@�����*� Ȁ��'6
96hק��-hr���"Q�c�~JF�ہ|��QjDV�n`*e�I��>+�� .%`F�c���6D	��ڃt��%>=ʚw+���Qe͠t-@���E����̿^��(D��"D��q[`��8�h��$O3'H�*����`b:�A;1�5q (��&@x�H��KA�����!�e�Z.��<�@�i��i�j��dCtI�a���^��I�l$�C�,5T��m��h�>)s��S�O��[�a��o��|.|��g]@Tn9I�� �;zF����å\q��@����g)���=j@�V�H����Y!�I��"*WD\�&o䅹ChN_≨8�N�H��ɮZL
 �"�@������@8l���Y�%�" �����
d�frrP���1k
��[�h�|Z@!a$#E̓\�� "�/�+����(ș	��ʡ	"&�ZͣB끾J��`�����>O驐��(&�@*'�ЈOܴ�C�#�P]%�ɏ6���cs
JU�6��K`D0�׎�<�N@�ǫZ6���E|"@�%|���:�O_�w��՚TE�%�TYD|���1��U�zӪ�'��׍^�=W�1<���G虁<]���w�'���;98
�R�ڔ�`���I �b�h�>�З	d�n�ŅOӴ��U(��a�����mX��5�2ƅ*j>��ːV���im�+T}�7H�Q��1��Z�^�L���+k]pW�F�1O�U�^;cȪt�qń�PH������?�#Z#Q��Cb#X�$`&��E�	.dưeK�D�K{`Ei ��"Ȍb�D����=wr1.ĸ�%,x����]��0�3�8"��!_�]\�pG{D_�wh4Ҩ	(k.t`����+���yc�V3`�����2�p�V]��b	E}�k�f�ڕ be -6ґ�֪�$_;�`k"�M)b��|Zc'�����&��0��]�.��1+�}R�üE�ʜ����I�S��tJO��fl�*�HO'�r�p�HeX�� Q �����b�,�
��z�N�V�>lYW��<9�搰p�n�h�DP�ʵ��iۚbE�d���	u��&g��
c푾Eض�v'�86���$Q�pV�dK!/�2�awa�'�D���'��x��ϐ�B�	2�	��OY�}��4o]x�Q$��<���!ۙo�R���:��ٲ��<BZ(`�WA������hyy��N%!�x�$��@C�j�V;���{0��Z5|T�t��k��!��GC��	ϓE���%��OWJ|�K�/,T�x��Y�0Cß>�R��9�|`��O#i�a�O~�ɚ!9�g&�,Inֵ��R�lr�tHT�I�zJ��1U�TȓE޳����Vꨫ��94)� 9b���!�ȱKb�'�>�A���>�B�E"k��T�'���#tg��@+�ٱ
Q�|YuQ�@��%�TM	����۷�	I	U�AE� Kl�� ��
)X����?����I <�/5Мj��8�B�Ha�_?(g:is`L�#��X)�o8��
�;����@O�1�L�"ݓ&#����x��u��I�g�F};�	��U�S���.�)D�ђj��\�T�.�ɞo�z���^��\P��eUJ���׿�?15HC��v	�%b^�l�L�'����cb��~����CԜ0Y�!*O�5���*L/T�"�E�}�>mZe�O1gl���J��ir^��S�Æ���u�J�'�RT��̈I�0�ŀ
�~�;''U5h����� Ӟ;����懚��d�Hs�b��7'�-P2Q����:Ny:�P�-��:�� 1)ux�X�$�]����Cb��v�n	J�.��r�5K���O(a+��<a���nM�{��#� ���	YL�tlX4��m8�|еi�<7��	�v~j�Bm��-Jĸ�Vg 8%�	j~�g:-�FP�hئL��+��q�
�6���D���B�jU�FT���'���+��ŊF��	����1=Ab�� ��\d3�n��hES �=}bl�"��Ј��=��&J����'^���Wk�z4��&8��I+O����@޺,``I9�/ݿ�����I�b��͂Ш��'�a�@��rb+��HJ8�uJ,��i��'|��b�T8aX}
cM_$c����`L���Ї����Ovh���kY�(R�7m��["iZ�a��L6���d�����I��K� �pp����>@p0��"�Q`� p0�%����GXӺ��O��qnE�35���獏��D���N~�'�
��%�/��mb#��.6z����qX�!��PX�5XQ�ݵ8��O��+0�Y�+���B`+�hU�?!`�Q<V'V��H-C��Yqǣ�7h��m�Oh��ǚ^ݾ@!�f�S���i�g��{�0yG@�-u�\q��[�y�X	 #}b�*��e��!$䆚.8���@���?|��jIDC~�p��܍O�������.�㟢|��ǫ8q�lk�AU� /�aq�(�z��/ޖ�T���+���N�
}��`��'�.I$8E�1��x���<;t� �J���5E�IR��أ���@�:$Zr� �I�2L��Mn�d��B���A��ϖ! ��i��\���<A��߶a���k��L���p�'��&��:�o�I
̩����BR(��dJ�sy&��Ȍ*om�q��ə�D���螓Ʃ�mL�<���Oƨ�e\�|��+�C�<<�8���$F�5����ǝ;{��T�S�R<	be��]�н���L��2�入t����+��%b�%�	�^����4!�	�{�? *���%DǢ�)�)
 H|�1O�h���Ȓ 1��쁗7���b�)�I�"�{�I�c�A:��ϓG��'L�t�s�O�*�P8��슲F"
e�
ϓjAP9��䚒�
d���Z'|�r���+$�܂��c��W�\}8E����h7�<�\���'ڸ�$nŝ.����оZ(�BI<�%Ɓ=��Q�J7Ĭ���B�rԬ�"�H�'�X�[bA˞2�M(���*}r���W딽2�bQ�{�����(Lc�Xy	ϓG����������R�|����)����pCN3��;��6��`�:ݒ�Ȝ�i�TrR�@V螩�Ī���xQ	bX\�Ԃ�Y�C�X�y��OZu$�� -A}66=�v]e�hB�+�	;�<a9�IJ�ZzlmxD��d���'�
Y+ӄ�u����b-ӎc�V�B6���r��[c@�lV�a5�I�]G�	V��KTﮉIS���$S^�bѸi	J9�D��q�갲�l:Ol�`�o?d<�*������j�wZX�OT���Q�$�ve�q�b�/x�q��8�(Ac�G�x�s���y�c`6"���W9D,�+c��Z��Oʙ��Ǝ)؀�'���'^D��#0�J@�Q�T�6t����Ƥj���@���;���#���B)ll�&˛ b�L��S�i�:��f�,""��1�ۤ>:ęJ��qǛ���d+��v0���'*P�ǥ��C�d E%BGb��p��<���x�i_$�"�sP)֊I�*Q�í����e�=Q�CȊ~��`!�d�%�8�Pΐ���D�LpB%���0<!F�� �`�q!�كH� axqM�+"4X�	`WZ���3C�`��ꊔ�y��qDhZ2�e^����BQ/h�Y�퉒vB	�Ab�[��_�o���%ƣ`��q���;�n��Fe�x[�'[�A�Sz����H���)`�W�7	b�Dz�Kǋ-��})v,/����ڻD1d���Í�\��hB�Y7{V�s+Ԃ�Z��a%N�ft�ds�oE0R
Š�x��R�' 躜�,җ����7K��y5�t$���3C��9��u��ۙaH"|+�b)�i�F�{�����P�ʗ����҂eվ��'jdI����O�Y(s�\�B�Q�gN�[Y�}������l߼n7�A��EGK�nu����Oq�J,�c �?n�Z�!�GJy�'�أ���cX�4�B�*�t��/MWc�� SfV#o�La�&E�.z��dY-r�f����3�nX/���Z�IT�[wM�D�lױ#!��,U��0�T/I6:�,h�"N 4,��3Ou�e��ĒhB�B�J�?���>QpV?M��"6lA(�YR�J% ͸��;O��oYk,a�0��+/�2�
uG�d�T� 6�^)�h¢��3�pC�I���5���!H�*Ps%�;Q+�C䉫F٪��O�0>��XBFҴͶC䉑}��K��ճN�z��Ŋ͏y3\B�	1v���0�R�D/D�pp�E�S�&B�3N�Z���I�6�Q^&uB�;/�H�{�N�I�2�T:KBB�I HNF���v��mӨ[{(B䉞 L�x��+�p�e�D(�:�TB䉝>�4M:#"�!f�$�t��� �(B��JŢP-������f��7D�@���.G��ŉ�'X��A��k.D�|����?�"���9v]pC :D��{"J�&zR\�A�B,G6Ek�J,D�Lwb+@T�E''g	v���b(D��ɄjNC�PD)��B�{\���8D�Ԙ�"/̵a���YN8��8D��)2��)dF<��E��w&6x�!D��Q��_$
��xi�Q���(g`=D��*����˾H��YRCI'D��(e���9�Tу*I{���9��$D��I��T��U��%M�y[(Q�l D�,+r.�3g�����IP�c��a
>D�4�d���N��"�EOq�����6D��1��d9~�h�z�Xs�N1D�𫵅��rn�̘�&E(N�R�)��"D�Da���B��ju�X�*4�	1ք"D�����@��E���I�7"CҢ%D�L��O b�(���a�4��eʷ�$D��x�h���a'@ذY����#D��{�I\�E>�܂���3h��;a�?D��Sa\�+�z���`T��Xi� 9D�� b�[�i�&q:���
�L]֌"B"O��:���x��(��ԗw����"O⥙@P��Щ���
8p�9�R"OqRdA���l�rWf�;T
1�"O.@���J�pa�X	s#��\<�ų"O0}0��!�blC�`�1 �9jB"Ol���2K��iE�/daPL�v"O�H��J�<eZb�zf ~-�Q#"O����C]�h���]&9�p"O������6���U���% ���6"OH`#G���g���tlHj���V"O���$L�V,��b�Hj����p"Oj�'�0\���;sI�+@ᣂ"O�2�&x�d8�E)T5Ґ�T"Orq�P-]�j0��Jǈ!r��&"O�I˔Á��"�q�Hնb� ]�P"Oh�ڔMH�?�qQ'�0���"O̱r&E�"�p6AM52q�y��"O�XS��+X�B��K����r"O�$hwDY�>��YI��Y�H�f=I�"Of� p		�w�N���R�Xu�Ab�"O�0{����.����C����"O���k�N�4����L���B"O�]B��>*�h]�%�)lP\��s"O� �I�8w�������M
�"O$�R�\�7��e�7�P\���r%"OU�C�W�a+w$�8I�(1�"Oxb�C�$2��q	��H��}`"OBt�������+�,)9��.D��@�ނ.��ڳo^2�¥:��*D�HB1��W�jŨ���\ߠe���3D�@�F���<@@BX�e��0iS%1D��A�H�.����f"V�f��,[�n0D�����(+H�r�S%sK��@�(D���qʒV�ha�O�6���c(D�"��ǍI���ó$MSx��
�<D�8�V�NV�n�+Bc̣����m9D��#�Nޒdy&0(WE@*��#�,6D�,R�ߦ 
��є�U����s(=��0<��㉕7s��� �,���#�BL�<���]&R!qn@ }|(� ��yB��%T��ha�E�p\r)�1���yrg;[R��@jJ�ey@dP� �!�y�i8��c�71Rd�����y2���NFx�+��*�v4kE �6�y�j�7�hI�u�/.�+���y���jp�aG:mt{� ��y���:܊p1������*��#�y��N�S��ԉ'.�&c��U�al���y�-T8c�24�Fޘ-I0੶�؀�yb��Iefi�&�<�P��5K��ē�hO���+��ڡ: �g��<B�(�"O2E�vG�:*��9A�L
?�$UH"Ot4f�Rl�>�Q�A��"V�4�E"O��+�;{��Aӡ��E�:r"O���#��O\l�v�S�bЎ�(��x�)���*$��#�A=�&h��9=CC��!-r�yQ�ɳJ��5��R�z��C�	�Bjf��C�T�1��� �"z,�C�	bC^h�7h�"a� p	`��w�C�01�� 0IG������-hxC�	�0�YS�DN�5-̥ం5BC�	?Hy�ӄ�� c�]�e
I�~UC�I87�P�u������J�-n<C�)� xT��J@���Qڷ���9;��I�"OD�Z�b�r��@
��Q52H� "O��J�/ =��e�2	�s3 ј!"O�T���S&��g�/���p"O,�2��:��T��&�@րA��"O��sPn���0+%���"O�a����R�@�[b \5`�X���"O8���		#TUS�R"�̀�"O�@&�ĜIW�pW�Y�G�ڴ��"O�(���eG��Q���NR�"O k��K�Ofj��AA�L!�"OJ�k��ƈ�8���)(�t�Hb"ON�YQh_�&��[��]�T���k�"Oh�RPO@�=N��x@b�lW� i�"O\1I��N�(�d�1� ܫ�r�r�"O�yq�E��c���b
@9@lz�"O:H�7^�^X}��&f��h��"Od-�L�zSD�'���$��hr�"O�|��K��=�ܳ��\�r����#"OVej�Ɨ�^㌰�q┯B���S�"Oڡ2���	���WL��kۀS3"O��Rb�@r}i�ʌ��~�ɰ"O<��aZ�*���c���Jc"OX4Q�C,_n�臊��x�ι�G"O�����(z!&�[*�+��4;�"O�$P�+ۂ5��x��	�
���"O�d��ͪwOD	��˰v��t�Q"O�`�d�'vB�̀צ��?Z\�
�"O@H��%'0vd�s�_plB�!@"O�5!�X�K��T��Â�C����"O����	�Is4�#q-H�Z�\@H"O� �J<� @��a��xyF(��"Oh���l�+G��q�B��Wb����"O����\�R��E��4d4$�"O�s�C/`���Y�hZ��A"O�s�R�M(�9�0��<Jr�A�"O>D�E��:Ch4�#�ܓ����"O�i�r���EOb\��A�l��[�"O�H��8fQ	�!����"OL+��ũ3L��ҕ�T�S&%@t"O�9����a#�I"�E�:IP$1"O.���#D�;�@���d�\ό���"Onщ��٧H����Հ�,,ɮ�"OJ�G�5��!ڷ�B��
�"O0�XFf�<<��O�;8��'"O�	�D�(d[h���@H�#1"O�跪F�"vT�"� ���K�"O�p�Ղ�4�� ��k���[Q"OD�K�f��Ԇ�І˅�Tx!�"O���,ٺ��;�ib���"O�p�[h��o���^�(�ȏ`\!��	�(t��&դ�ְ#�PKE!�d��~L����Ϛ�k����*�M!�O�d3�S+\�r���|�!�d@R�"�C�C����bϓs!�Dt|Ab���('�JXJ�$
c!�$�e����J
=^ޜ8�e"J�e]�ϰ>i��հx�1��8����j�S�<y�#��nɺ�e�
%q.�e�F�<qF��wLai�k�]`�����C�<�V�]�g? �SQt�(�����H�<��-�Z7
�k��"΂!1C�O�<a�B��,-BH�4i�9>�@��R�<qB D�?��DA!o�y�H�`N�F�<� "@�����eM��� X��R��'��O����O�	6Iք �L��d"r"O�#AK�pY:49BFި�ar'"O�4���Ѓ5|��㥦Ϋ.��"OR��AO�_�ܵ�%
5%>h)�S"O�l�%��{��´�Z:X�s�"Oҹs7�?ʦ��$>��Y�"OD=�HZ�I۸��b)S�H�,��'1qO��舍�2�ӎ��8�*���"O�Xq�4w�,u�*Ym4���"Oh�i�`E��:�IC�%i�P��"O6�653���n$/�%���&�yrjW�Z����w��4�#A��y�f�<�艸�g�+v�Mȃ@���y���e0�S�M�;��"s��,��=��y��a�<��&�#8K�M�(��y��>k�TZ�H�>�@�����HO>�=�O�,��A%�<W}�=a�.�0�\��'�L�b�'�2�6}��!
�&ꆁ;N>�
�G��p��d��=t�w*�n���GE
}A �3;���*�����%�41IGɩk��p���o^\!�'/ў"}�l]�:a�v��X�4<��@LJ�<1�@�.8	xi��b�2�ƹcTq�<7�F<|S���)
��A�u�<Q�*��"��ŋ1��
-, MD�As�<E	�� A`�K�]D6Uh�hD�<y�KY=`k^U(�(&-Z|��DKt�'6ў�'c� $A�d�x���kE�z���ȓ~'�`����Q6��t���2��Q�ȓ4��H�o�YB��mgX��ȓA�|�Yv��#��1���U�S���UI������1\����`�	]�ل�l����X[��P���4E*��ȓ4��#e�=`��J�	#�ȓy�H0s�!eU<Q���FP���`�(��PF�Eʽ�%j�(��чȓ'�X�rq����B;�eD�"��x�ȓ9-���' !&x��"0��>B�a�ȓ@��	P[Yިq�6��[�&Mie"O�A)�|紁�KӤ|���&"O��JT��,�:�8�kQ(>��x �"O�X)r�ظ�
�R�����ڰ"OXP �EP^Sɢ��z�8xS"OD�)�JF�Kf�kB�nn��"OrTx��}�*1ꎌcs.u� "O�P�*y ���)X�T]LsC"O6<�u�̹ �H�ƛ�:PD��"Oܵ�`写�L���o
�H�!�"O
L� �_fȌ�<H(���"OX�I �֨p���Zl� $ߴr!"O����-'8� ��A���PYy�"O*H:��]
I� *�N�6�.Ԃ�"Op�����8`���p��\t� ���"O^��2OU�)��0����|pK"O~ 	סĤ/&���uC�vd�@a"O2����>x�I��O/q_е3"ODA	��V���!:��
V�|;�"O�xcI��+�&-�ff�0Bl����"O��Zn�`����ę!r� M�B"O؁V���qva�#����U��"O�Id��e�A#"�˖1����"O�H���7|���f��#r�؈"OZ4��J�� �D���.ey��*�"O� XMR�6}�Yit횩iY�+W"O�"L�Q�.�J�A��ve�q�S"O��ҕ�R�(��h��K�VHHT	�"O���K?C�}�@�"I8�P*O��+�)�:v2��t��#�^��'��/^!G Y�d"�k���'�(* 	�LK�eӠl |t�
�'kT�� �(���Be@Az��b	�'W��r H	JW���%.�KԞ���' �y��G�'f� (��[�X:J��	�';05�!�.=~�#6ˋ�F���	�'f|p� y~��a!�1�")�	�'Z�U�Z�{�n��4�ŝ����'��`@Ɓ�%�`��A,d͑
�'mȭ�d��;͚�`���.5`2XX
�'�p�BG���Ґ��b��+���z�'@��H�+��Y!���<we4A��'��RTD�-mC����L)m�B��'|�DБ9*�@,� ��'cn���'���2���4hT1p��$M���:
�'��1�ש	If�9ׯ܃6�A{	�'�Ƭ�B�ԚEc.P�6�� ��$��'�`��"j�H�4蔔jL���'ːY�"��0;���	T�]*l��'Z�94�&vZF���Eӂ �F���'����2�+F.��J���5} �8Z�'�<ٷ��Q�Q�m���i�'T�cJ6[�<0àL8s�|!�
�'�,��&�d�ȵ����3:����	�'R��RP���V*J��qB)(�x�h	�'=��jDc�ZƠ�o�%W*��'Lpp!�ߥ
̨P0�kG6l���'�R̉��Q�pn1�҉l;&H�'CR�������g�@hb���	�'�d��a�m��aH2��;b�lJ	�'Y
-@�!ޡg0�a����-��'Ȕ3#�Փi�6�x�H./�\�'���w�6.������9��
�'���Q�Ԃ%������@-�=��'��,�!���G3��+d؀1��'�J�!EN�-`��h��YhI1
�'���!��/����ȘR�2���' - ��d	�
%�E�{�<�B�\��h���)�t�<�,�w���7qlB��E�Kn�<Yƭ� �@����ۍSǤ�¥�a�<��߁t�r�qgH���keKe�<٣*L��v�*T���yB��a�<Q���.t�®���zj�e�g�<ɣcvY��2�����6�_�<��#�.0Z����7~��L�"��@�<Y�p7R����g��� �{�<1L�@R>�2bN��I(�XpЌM�<9��F,?�L�3�W�$MvPh�nO^�<ɗ+V�y�l�f�]vL�ݻG��V�<�1�8h�,��r�ڈJ4Hi�d�Tj�<�u&W�5��k�̏00~$3�f�<qd�L�0�bv
	�O=@K�G`�<�5E-]�X��K@�d��=�h^s�<٦��.H(ՓֆŹm���$�^k�<1w)D�;NR4 �5RlŠb��j�<�'�ЪN��!�%�/t=����"Vj�<��I8=��x���']@�˳@Fi�<�SZ�	@���ܸY���0�h�<� �+"��)/"����غF��h�"O*MѤB�:�z��2�
� �8�@A"O&���#�0~���$ٯ%�ތ9�"O��'Ȋ�	�r�+����#"O���e��v=Di���ϪC����"O(pN�e�JQ�!�c��AH�"Or\�1�"��� `A$��H[�"O����dϵM��}�`�U!�x�ys"O
�J�㛑o�v�����s��}�f"O<ű7!_9e��ّ�F�.��`$"O��)��;��$��2Y#�p�"O0��c^�B�r���-���"O�Q�&/�&�p$a��2	R��"O�x�іQ�� +ՅS)XK��K$"O��:4����V�xA��8T"OP S�e�x�8=�0a�0N�a`"OJ�*T�[F=�pkկD�b�BY��"O��p�ʟmNH��)[+�@�[@"O<�����x, 6�	?'o�p�"O6eJ����F�03GT�/\��c"O�M(�Ş�g��uIp�1���e"O��+�#�1Cg�LX'�Ӝ+ޜ�p"O����[9?�
�1b�>&��"O2� �|:&)1�@�n��<s�"Od���K�X�딮�"��x��"O��ʑ��|2ܪ ֈ�Fy�S"OH���灷/%��(���p1�"O&U�^!'���!��^�^���"O�H�0��p��p�7�c��5�a"O�l�V�<`����wK B�Ɲa�"O`y�M�4&K*ڡi֐���"O����F3_ �}qe�U�CZ̐c�"O��Q�b�p8��@�'�nP�Ͳ�"O��0*�ܶpVf	�4%�ԉW"O�ԡvܜ�
� E:��(6"O����,�,w���.�x0k�ɏL�!��P�z�� *7/%I(WI���!�d�:v�z��FL$���hJ2�!�d_wFk�GX�J��ErC�Ud!��E�t� :q��.� <( %]l!���?*q�� �·A�&�P���8\!�df�@�pF
L7ktT[��5(�!��I;Fy�tx��^+p����Ӽn�!��:�H�-��N��}�mǾ-�!�dK�'=�!bKH/x��@f�%�!�q�zTТ�'b�deh�&ǴOS!�O-c�];�쁹f��Q���w!��)9��a����/��E�׆ I!���?F�J�3���1�$+��W1�!�DϔE�`#%��.�%Uǝ�t�!���v��`�������څ�ީz�!��?��dK��H�m�D���!��p�^��Vk�Yc�aJ"_f>!��Ѻx�d���մl�܌��S"!�䍞	<��f����`�`ՠ�!�$ѵv�\I
��A9\8<�yef�0�!�dH�T��9� �ɘz" ��f�9E�!�d $5����J�!��H��!�$O�q�i�#�ؠ{����F�_=!�dH,R�"ْ�C2j��!s�b�ў\��Ue���r�^�~����� YL�B�I�5�>i`п7��LZ6�� 5r�C䉊'PZ�H��"�貲oW~��C�ɿk� ���:Mݲ̡@MW'*��B�)� &,�dM�'(*�"$�}�|�IE"O��V�ؼ;�в�B� �@P�Q"O8�Y��F}:�Eҋf�X)+A"O����k�W.Ը`!o�b�.9�"O��"��N)t�"T��.˙e�bC7�'���,B�L 7 ����3j
5S7!�$��ܴI3	Of�V9�*��q!�DZ3�"	`�.�5��4��� ^!�" "�Y����j~^�A�Jݚzk!�$	Jv�:�I5}�)� �acџ�E��k �A�Y�%@�:�B�+[��ybCA�qg*<���� /��ڗN��?A���Ӹ$����4��)���A�μ��)�ȓyj9xrb�3GW���' ;��݅���X�4c {I� ��� m��}8���2��)IBG#V��ņȓA�PL��� H4j�CHQ*"�?����0|R$�H<�(d굢�
��h[ğv���0=6�*pR��B�%j��C3�P{y�|r�`�ѕb����Qi�=Q�!0�g5D��Z�y�F$��+�*�xz a3D�d ���+:%h�I�n+�1JBO5D��ʃ@����p��Z�7�dA�!�D�gF>qcaNȠU����v*]!h!��v�E�`�?y�\ԑ`oG�A��ן�Ih�����OP��By��난C/iWi�Oj�=E�$H 5 ��b�U�H5���V�#U!��ź; �!.s�T	���A!�d�gk	rq`�kĴ��v�ڵ!��e��Ua
��0c���.w�!�μ�Ҹy֩ՅmOtA �M߯�!�$G�_|I!4LZ�?e�%�7lN�v�!򄂌Q�nEqȌ�x��;���!�D��9�Q� /�LP�f��f}!�D�
�1S����k耪��*q!򤉤#�.A�N��.�X��L�q9!��Eg�`���NL�:�1��М7�!��īl�����ݔ@� 
I�V�!��N9b����g�@iu�
?!�C�w<�����\�v<�L�d/!��Ƚ�j]��,]�en�{Šȩn!���rbԃGl?X��H���=9�!�Ė�z�j�~�^���W�!򤅈Av�Q[wG_;yP�#�k�lr!��S��dmx�i�"�QT�*!򄛺V�"`�f�8|���;����!�d�+mVޑ���N���:el�J�!�$ݯ4}L�c`�0����+ҍg�!��X�@ƼBG������X�8Xa�'�&5�qa�7��yA�)#�:x��'�E��m�g�V(��$:Dƪ�X��mٳvM�)�(��(Å&ֈ����=�J�\�c�����v�J��6y�H��qV��{��� ��
�cQ.p����j�ǂ�5g��t���7T�Ą�cvdd�ł�Zy�聀���1n�|�ȓ���q4�W1Y
S��rp����p��ѧJ�C�= �H�8n؇�f�� �U��;-��!� �9I̢u��G~��#��!�H0B�B!�X��ȓkE:!g�L#E  �ň�9�̅�!�usŃ�9~�;�d��ԩ�ȓp���i���%(L��n�2(:��ȓ2z<��������e�`ń�S�? �HS�
�#�H�����	LR�Bg"O��#p��;t��Á#�(OI�U�2"O���M���w���$;�K�"O��9Ԯ�@���*9 0�v"O�e;�eH]4!�I�|V�Yc"O�9c�/dU��*v�[�M��R�"Ot�(e&٧��}�_')���"O���b��B`�G��/#�:��r"O<�!��,( 4
��p����"O�̱�-��L�xU� �M�h���"Oɲ� ����3�Ka�.��"OZH g*@g�;ԅN�.0"�"O,���	Dsd�_�#���:b"OSdBܼ/�RQ��hW�
-�m��"O���eˁ<p2!P��$~h���"OD)�%��&����_�6KM�"OP�p� "�rW6m7X�a"On��H��>��;W'$''��*F"O� Ҕ��?H,�f�!5�}�S�'1O�]jG@K 'r@!
3e �i`��"O�uCsB�\�A�"cW�=.vi�"OT��j�;�vl�f�H�8(B#a"O�!QT�Ja5$�x�	�G6��"O��!"$���+v�G�("!A"O��* ���4�  ņ%	���"OP5��GF��RĩF3��U�q"O1
��`Z�	"��G�Z�|8�"O����.iN��g�܇���	7"O�XAB��	$ ��4�)Q~!E"Or�b�m�9M�ٰD���aC�"O:-Pѣ�'_H.����ɷj�u"O�q+G�� ��a����x�!1�"O�������T)��bŴ�4i��"O|��'�0o�4�c�M&\� ��"O԰T+�g��i�Aa��6rŃ0"O0�rqFɈl$ �J+0��d�G"OҐ�`_�k"@AR6O�$R�u� "O>��w�Y�dڨ����T�h!�K�"OL� ʀ�I����+ �s�Q�"O~�#Uϙ�!�<��PA֘��"O�Eфܚe�T�3@T�(y�&"O�q3&n�'F�P��O2i��T�"O����ᓾI"���r�P)ҶT��"OPX�JA_�f�@UM2Q�����"O��v��Y�萃��JyS`iC"OB��<�mA��˧;"	#6�	|�'��D%Z0"��paׇC-��"��B=e6��r�����$�(�ϲ&������V/C�jB�	�.h�CǗ-^t�+Ult�|B�I3kh�@���TT��C*�	v dB�I�c�(��׳LHTdRA���BB�	+"e�8F��_b=��dK�'g�C�I�[�p�2��[�C�"͠�Ǜ�-�B��*�NH�E#סp����ה#��B�#:�}��� +������܊B�IQK\-6䎽���3S��6D��C��?=4�I@ޘ\�|�h�Iٟ0��C��?F��С�l�$ր0��ʺu�pC�I�7��0�5zg�{t蝷Z�VC��Jh��2m�=e��Pԭ\�@�HC�I�q�z���� �N2� �,C�I/DH��߻4�(@i��J�0C�	3b{�����Y�� Q&z!��


�JQ�Q�N�P���B��!�� 
��%�@�NF2�Ѥ �$���Z`"OHj���,B$�L�;����"O�y9��1��=J'i��v"�EJ�"O�y*���{(����� �����'��	�iX�H ����uHZ�**�B�I�_��HCs��m�R�� "�t�rB�	�?#��[q��.]�JЀ!�KS��B�ɧi8�!�E�)/,��+�mrC�I�+��Ic�'łqD����AZ�B�ɥ��a�F� &U#T��(�/�B�	)d)l�G#̀O�F����>����O<�d׀�+/�8g�>(Eb�->��A��;TJ4��M�O8T��,,Յ�� 8h�b/W�
 -�*qޔ��iJ 4��\�3ҸX{�J(|���ȓ3�1��`� $ x2f%ώi�(1�ȓD�*�Q�л&��2CQ4l�H1�ȓY0�;��OT�BY�ю�tJ��G{��3�h@ �!u�"A�`L�4�x�<y(���I�mX,���u��q�<P�_�=P�ESB��s�>���'�X�<�P	��P$�lyT��>�y��p�<a�0@�����BO�vh���Rp�<Bm��&"�gg�G�$[r�S�<qDJ�e.�((��B?o)�����U�<�`�	X�T�b η]����iO�<�U䒀n=��J<I�� �Ы`�<ɒ�H� кQ�Z�q���^�<����\d��A���Lg��	P*�]�<A	3u�����Q�)�2@)r�X\�<�P�ϓv V9��:!	�q�R/�T�<��� k��a #h��F�r-k�)TM�<���=:&��"�)œ(��$[��T˟��I̟0��	���a��4b���Ц#ٕLxrB䉩+���"��E	-��6�{A�B�I6\���NX�>�|���%�=
H�C�>v��	�6�F�O(���@���B䉽V�R�B@����YN���B䉟��d�A�!����+L��0	�'�0 "�ΐ��Rc,Y85�y����=�OpH�"���+�.���?zD�4"O��:��W�[�Xа�R1	)�%+�"O���L����h@4b"�U@U"O>��q$͔C�@8��a9Jl �"O�qYT%X" v������QR�'"O`�ˠ#!���J�`��Ј�"O��KFM�W����*ͼ�bG�'R��'�a|�Z4_g�@!Ԃ�%lA�U�R��yOE�T�d2���a$�\��m@�y�B .��x���>G�������y��J^U��b�gV���0��!yk�B�	�
9�qyF�@=RhzlIV�V1"	�B�I�M`�x*��� e�N$R5��3\L�=I�'B�`$�5d
� �X�C���f�Fą�J����@͆�[���v/��Y��<��`�&Q�@���D ߖ0k���ȓd8)@0���5���i�EB�NW�e���4��e�~�yҖoŁE����ȓvL���
�"y��	�(гޮŇ��	�3�E`du�U.Rp,�ȓp	�x�ҡˌB���I�1[�Շ�[��C��'Ú�P�hO�ߠ�ȓvH�&,�zX�H�Ɇ!&:]�ȓHȬ��&���*P����߱{��)��S�? Y�H̺|64�	r(��C�����"O���%�WV�D�����Q"Od��c(��R��C��4��U"O6�w�SC��lSOT,cŠ�c�"Of�Rb&� �>1���>���@"Ot �хS�r�8�V/O�a����G"Ol8:4fK�g�%AS�^�7��a["O89��*�	�R���Y/ �a�"O�����?y�W���<�ru"OB�A%j|�
a )#�,|H�"Ot��ǒT
ěD��!�8���"O��Yǃ�Ug��B�� kЄ�["O�\9pȪ>(��P�h�E��]�"O�5���]<C�`{�]'uD�XKF"O�`S&�Ǜ���T�K_4p�J�"O�I��
�?�H	�� P R��"Of��da��I��̈���X�������$��ʳ-,�Ԓ`�#�
%˳i	X^!�d� 0�&��N���	f	��[T!�$�&�����@��f@"��މ0R!�D��+挙
��	W���k#d2@!�"t+n�.Ƹ���/5�!�d��Bj������&�,pSJ)D�!�$V�	�3e�t�X�:�!�&	Y1O�5�d�'�Dy�"I��8���.0�qy
�'�D,�`$�7F��P���	�"8�	�'j��s��&,6�x+�yeLlK	�'�ve����)	�`FJ�}�tj�'�l������$�#�a�xFZ���'��!�Ն��I�6����lZ� ��'�8��C�U�R�����o�S�`D�
�'#*�����M���Ӏ%��<y
�'&ލ[r���j�+F�.b���	�'ͨ817f��cN���$�A]�p�y���6E9�����K�R���+�y�)�5g��4�'"?�<0�KQ(�y"g�*I��X�UdߐB>xPґD*�y���Z��E2�cٸ8�YpN(�yr�i��1�C�{�h�g-�;�yR��0�Œ��U
,Ƚ�1��$�y2�	>3�8���YXfy�3M���y�fƼd,�u�,
8~�d���:�y�@^��X�N��t�X�R�k��y�iƐ!%�Bb�%]�,͈r���Py͟	X�V�rr)V�7�z�x�^~�<Iv ��)����mD~]J���~�<y@��6��qe����}pF*TD�<��نix��#%V=J�ڃ�G}�<��i۳?CZ��3.�iZH����r�<�F�Q'Z�д�ڻȰ��G�KC�<qu�����/`I����g�G�<�aH�!b�P��P�C!F�J�+��C�<�S��09��q����D���ǥRy�<���O	D5��z�k�j/vqKD�Ix�<�'��P(�ƒ,�(��P��i�<�1�1
H��j�F^��c"�Kc�<Y�e"Sv�X�⇝W\$�`�[�<�fB,*W�Y�$�m頽�d&W|�<�VID!��# LF�d��u�M�<Q%��D^$�7NV�W���;�lDQ�<��G�~�|�
��0�$*�BG�<a�,�C'D㱆�*'i*3IJ�<9W-��"��e�����"�LH�<�mϜRQ�@0d���&BE(�LH�<� �j��/0��c�N�v�\�˒"O�з�H�=�$��rmU:�P�`"O(5H0c	���)q@�7D�t:"On�pF,�(40�W�ҢF�șd"OzaIE���\;$���^!`�2ls@"Ov�ECD�lN:��J��P�� k�"O���'��+�t����ˎ$��M�2"OꌙAN�A5�����H'*H9�"O6�:3,ѕv�V4ğ W�$P��"O|�#���;}!.@1f��8�\��"O�m�&E,:�d��J}mPAȔ"O��P�j�	4���)򪐲|a�xh�"O
	[��K=x���!i�(K��	�"O�VS#fkfQ������ySn�I�<��mH�_��낧�1�:��B�
a�<aeʈe�Pٗ�E�e蒍���g�<��$��-J��Ʀ�o�0��A�}�<15�P��~�q� $mC��^�<A��w�������;g<�:V�U�<��+�d��1z�$EBZƬ�%WI�<�vD��f�X��g�s*��`I��<�5.(Z�Cs�u$�uR�{�<�#pa�
�Z�T�"�g ԅ����Ƌ�y_^� &+L�O<��ȓu͂6L�./_�p@kx�T��O��`KOn�p|�u�I{3R��ȓjZ $�d�y=��P *��8��d��6�E����5m4�R�LVcx�L��i���cZ=|K�T��1W��Ѕȓ���_ l��qA�<�
�"O�e(�I��E����
�a�"O&�8r�N�(��q��fR�!�|U�Q"Oj�0��e����E��G���hq"O��N�.}C��x�H%�"O��ǜ�1PF�:6d�2tyJ�*Oऻ�JDn�"�bVi�_�&�x�'\)Z���F�h�൫ʽ\*`\��'I�d�#H��t�\h�(M�MI�u��'/���(ڭR��5�%d�#C�8
�'���*�G�&FqC�X�+����	�'����!�*$i�������*
�'W:TN�j��	S�� 3���';����T��ʽr%�C�H*���'-�da��ED��TnU�0��'!شC�,p �Ж�$=yt��	�'��%�f!�1+��IENM=5P
T��'�@�[�Đ�`b�D˃,K!��	�'���+��%A"9rc�#�	��'��{u#�<s\ؙ��B��s�6,J�'SR%�H�
<��܈�B�?�� �'�e���B��9�h�+,�*�'~���r덉ew"p�q�W�͠�J�'�<�����:`�cƏ7�|��'�r�+��� �qB�:^:V��'<���*�X�ህ�)��Q��'w\4�&��Bf�B����&}t���'��<QC�ܶw¶sW�Q<St���'/��@�צl0�ܰ�͍�j���'f� ��\h�.���: k�%��'���Rc�vj6�Y�CD5rN�Ū�')t�!fdυ5T���F-ߛc��$��'4�����
 �l�&Н_c���'/���!��j��a�A�W�F���'F�q�4O�p�� zP�Ϥ�����y
� J��L�lrV+�"��`���"O^�)@"H�:�}�'` i�΄Y"O��ƈ�f���O\�
�Te��"ONi�V��j�����L�h*ĴP"O@x�UG�)*��`�M�p��+�"O� �ƫ�]Tdl���Z�x5\�#�*O�����1�h%��n�
jT�K�'���r��
|Ͱ���#ժ��'�6�Sp�O��D�Gń�
�8���'h�q��g�]j�iB�e¨.r��'O���Q,Q�}D$u·CY� ��D��'�KC)}ʼ�@��ciػ �l�<q6��y���S�i� ���*[i�<�����Q_��R��*.L�
�c�<���� �N�##�&om��#��_�<���%YX\@@jݢVɮ�� _�<9��2����%$W�|��bqo�X�<9�&��[���P��Da:w�R�<��K�s
,5��)ځ6a�P�J�<ѣ� �p ��-�:~*��Pao�<	��N܅�
D9t��C�B�<A.���� �j�4*��nP{�<�"�L� ��U�R��/"����O�z�<���1�F�B/'1.�3���w�<9�%:
1�8�֩άi��
��DH�<����'���K�k&o&f�H�fC�<�����[Pe*��V*�� �FGB�<��M//M��ǝX~�`k�FYW�<gMT��zq�2#��"թRP�<!f�N���t���S�WI��⦃HU�<Y5��iӲ�1�1`�5���Q�<yI_8ΙR1�$ ���JTJ�<�A%�D� ����kg(<K��D�<�veP�pY�H�d �Mf̝�&FD�<��@�+Uݤ]��ƈ#2(5c��C@�<�!�>�u�4JO�~�6�:���{�<�T�C��|͊�'�'�QB�GN�<���ѐ&?�m(��χ(�X�A#�H�<�tME�ڕ�oτ�Hx��d$Q!��.���8 �.�ً�B��1P!��
Y�E rE��w�� =!��85&��q�L��@��@�'&�!�d�-t�r��ہ<�0I�n�}k!򄟟P̶�A'�*�&���,C�L!��ϭrn��Dj�#�J�����nF!��F�z�|�׃�o�&���j�i�!�ă(�fq�O�5MD
� ��9'!�L1=N90$`����k���'�������H����{ì���'�f��V�\-:����&�kxZ���'@�S���`!���w�(��'����R�\�]C��ѦT�j���' �Wk��V�T���ٍt�"���'�&���Q�(���V�P�i�6-��'S�QQ���X�;��4s�F%�'�x��E��&М�S�ɡp5�q��'��!����e�B����6-����'�Xd
S�E0e����r'͞*tT��'�h%	a� z���*�C��c¡a�'~Xyq⟖t�`�@(DJ�	�'>z����^cH�$
}��	�'ap1ۓ���|��$1�㕨 /�8��'ZnKV�Ҟ'�h��K�w�r؀�'V���$��l2w�
l������ �p�j, �Q.պm P�"Oޱ�Ԃ�=+�ĝP�-�.5Wl �5"O�a��B�|�H�)zgԤ@!"Om;���2l���a���4����c"O�!a�"�� Df���%rg"OJ�@厁*b�HQw�-w� Qӧ"O����K �"��c��k��d"O����ѦU5|�p�����9V"O|��x���b���9G"O��P%��@��%�tA�*0�d��F"OЅ�Ч\���mT���}�Τs"O�A��l�e�3��@�,�tAh�"O�L	�B>���D6�6$Z�"O�T�G.VCu؊��o�T��"O����
Ҽp��(����(aqP"O4H�g��W���B��JA"O���@��>-�����뀩%X>\@&"OP(z�� �Z�AI�{9���"O�$��hP� R�BC�}�(9�F"Op�p�[�2�|s$��*J��T+�"Oh�K���5ê����Ȧ>�rLI�"Of��C�n�0��!��b���p"O\���,N�0|)1��	��{"OAǂ�{�$�3E�D�X1zf"O��!��!o��X��[�� H�"O�=y*[�ĩ�Zb�h����y�3ƆUkWg� Q��B6Gפ�y�l�>Z�����Dr�E�:�y"� W`!)�C ���tf���y���r�`�:�O�(/|a�t�Ϫ�y�#�# � IsD�T/WT����N�y�7�pT���GE�4L˶k��yb�-	���òM�7|�P�E�Ӳ�yb�$`/�q�s-&c(�!�<�y"*R<}6����b�S����J,�yR�҉1�h0R7aL;N[�d�� �y�B.M�G�@�P�rP����y���4ư�`(�10
P�Sh�=�y��݉2�th�	�&����Lސ�ym@��rrdӡ"�N�8� Z��yrm�;��m��?���w�A��y�%H�G��d��h:���Bl���yR�
f�r��V�6��e�"N[�yb�&2�Z����/|C�A��y�LD�0#e2��P�X!�!I"h��yr�F�_/��q'b5R�R�(W*�y�Cԉk$��H�ÂRS��BU�y���!2���5�N�J�Ts��)�yRk�X(�ܸB�
0�H�����y���T�IgU2��+sG��yʆ�N��	 򢇓����&\��y���
0z��%H�-�����B�y��>6G��Վ��u� ���C�yb�2 �-&�P4gdи�hΞ�y��ǈd���*�#͋\#(5be��0�y2��F?N�)eOۀ"�d�$k��y�O��Y���߮�&�S��V��y��WiyB�ϑU8z�i)Ý�y���:��Y�s��z�����6�y�	��"`�e�6���)"l6�)�y����_Ȟ�`@	)��ugF��yB�P�8j�Ԓ (��|�d�D�y2���$���Z��������yr����SѮ_*	bx`��ު�y
� a���AK�J܉���(+��;b"O8@�O�Er0D�U
	[�>,�"O����1\�H��EF��P����"O*3!G؉>^�	s�@�#G�ĸ�"O����d�xS�9W�=|7:�P"OF�{Bf��I1�٠|�h�[�"O���4���7��cN�G�Pp��"O����V�m���R�]?}لi��"O��khŭRt�8dሏy���i�"O+&��? ���U�b����D"Ox�p ���H�|�9��q� Z�"O�tC��@�?���5
��#�H4�@"OЙ��
��̚�!L����E"O���$"X< �JM
$�h�q@"OʅV%د4�.H�6���X�
%JF"OZ���V�~{�����L�����"Op̀��}�t�I�$E;n���JP"O6�����L��X�c����V(�"OJF�Ŭg�mR�k�X���"Ol��$�Z�B�\��VM��4�Ԝ�'"OVm�@�9U�؉i�'!��q5"O�q!6U!f�bS-�=	(t�"O���#ǮN��"��ӁT�g"O��rt�ҥ�t��,�Y_4)E"OF4�b�GcJ9�_�"H6�P�ȓ[�����E���x�I�79)~Ć��p=��-EH4QHC��5Vд��W����"U]"��� �>�I��%z�sFP�f���PFK�b�l���A��Q��.H���{4�� Z�����s�v�RcO�7L!RQ3���g�P]�ȓ��MQ�$A�ICj��-�����RոĲ%f�
������
tA䑆ȓW|j0���?�č8��ʫ��X��^���X�
O c��3�O�6�=��ho���w͝��"���[�bԅȓ_Z����W� %cE�;..�ȓq��xaEK	:"�X�vgT��"�ȓ5��HŀٻZ�T��M4=Eȅ�	�N]	��ȝBX�ș@P�%ܨ��~L�i��a8���V�*S���ȓH�r5��9,d�pɡo��Pd��ȓC���p熏B�
E�#�ҏC�A�ȓ)2ܱ�ݢr�H
��Z��	�ȓ;��S�hp i��o[b��i�
)�	ZP\�H���� �8���23 !`C�1`x�#�?4����*Ŕ �.�	�$��Ve��1,��ȓ ��H!iց.��5��@I%	��ȓ\�R�A�$�TEB��ڢ�ȓu[`p3ݐ�ZfPEJ(̈́��K�� S,����ĄȓPF����鉰-��T���`�Z �ȓ��iC��H�CdD�ו�؄ȓz�`�T��g��I�B�W���ȓK*��8�J��}�*�k�ʖczjL�ȓ&	�e:ӈ�>@U4� k��Q�.̇ȓ����U�%�pH�G+نȓy��lX���C��@�7�I.��Ć�aC�$xfI�_-|{ É�Tz^��J��i2`-C%X�\\�EbY2H)Ą�ȓ�~�cS�ۆl��(e�P�:[�d��?BN�0�+�^:���Ȉ)���/a>�:6G	D��0�fF�>����S�? 8����J�!�()C���̼2u"O���T�
G�
���H1���"O ّ�L&g�`��FF?����"O � T��R-C��4.�Ju{6"Od�1$F"S{�yY��Ս7Τ����'���k�dM�h��a�NG+=��U��%/D���2^�9
Bo��gʤXZ#D�\:����Ly↍���pDsGo>D��ԍ�C|��.\�R��"�!�ǥl@���B̴A���u�!�ě�%�\m��D�f�v��D��,�!��$Z-��S��8e�*��`�E3!���Ǫ嘣��ti�\k�"�1�!�$B�*��	�q(�^g�����/!�D�8�]jǁ�/� *�  6z!���4[�0eI��V�D��]{��G�:y!�$��'���A#ّ{�t"��Q��!򄑷.:�Y"
�F|y%fQ�!�޳0��T�mV�5*�9)�e�,�!��~Թ��M�&<^����h�!�D��že����U��$�ѣ��!��I�\�4��D���K7��,5�!�$�=�T���O����#o� �!�䖥Y�l�r�ũ/��8I��b�!��ѷ~O�i�ҏ��#:z%x�H7@�!�D�[NlL��V�\HL �CX��!��J�sW�������{.�}PudP�!��B	�@P{7e�-lQ4��2/�!��A�a��wEH�`+�����*�!��b4�"�̠+�*`PY!!�$�e��@(�*�4F�<�֢�!���a����";7d|�����3!����W�qc�ȑ>#���"0aʐ\,!�$�!�P��*��|��q���	&,�!��H-8�i���8u�*M1���M�!�DO���Ɗ�<*�E
A��h�!��x�t���	?;@�yg-�E�!��6X?��*�k�3L�(��!��[�`p�1��'E�IY̔)N�!�?����V@�C����ۇ>�!�dC��B�rW� `�`��܄4!�p7�}��S%l���t���t�!�$R�A�~��f��&Ƥ(�LH�,.!�$��Yv�����Ȑn� Q��!�D�c�8x��
�-�H:�EA�"!�9=��PPcˆ7�ZP
 f�&!�Ę� �8C��³�~E��CY�B�!���`��qʅIϻ7���P��@�!�d[����RNۼG�����>|�!�$:.(�q��4�*4A�l�6_!�OG�8
G�ç,�(+a���V!��Y�iZ>}���� �2���돥�!���0�[�Y�(�r�O�]�!��c^ �(L$'��p�BcY@�!����6TRG��Z��H��!F-,~!���/x��Z"�ďc���xU��	-�!�䀩襫g�Ա9���"+
3C�!��+ Zb�OЧ�*�Zt
��P!�䞣v���"Ͻ;KX=x'h� k	!�D� 2p@|!` �hEX�{S&ء�!�DWiԌ�c��A�z1R	`��E�!��J�8L�ە
P�`/r|��΂��!���1@3D���(�^'h�S�̛�W&!�$S�tС���G� ~x`b�A6,�!�� �m@%�H�=G�[N^2���#"OPD�q')��${arZ�"O*xq��R?(�e��#{�4-	4"O���a
˟p��a��9Ja�"O���d��D8�Iy�i)�"O��֫F�`�M�$k�	U�˔"O��R�I1C�d8�	R�'����u"Oh�-�8��12�W(0�~urv"O�ј���e ����xaB�"O�EZwf$	4�aI�o
.�Խ*�"O���r'\��z�;e"e:�Xv"O,H�A�#p l��1�Λ�� w"O���`�;?j(�@�@
�ȡ�"OĽ����h�2u�CJ]=�jRQ"O��0A��,d����:�\�&"Ol�	s���4`�i��
]/�h��"O���`�M�
��k �S�#�"�#�"O���h�:D���1�O"��-+�"O�A�5��/��(rG��% h�"Ol ����	6k$�C��A�D�P�"OhEk� 6"�T�e+���F32"OtY���_i 4� d��v�T�X"O���f�rG�%��l�=)�鐦"O�xJF�C��&�B�
�#;�P��"O��g@��Yf�蛬��8B�"O�1;B���4���P�Z��*"O.�6/�4����+9�� !�"O���u�Qt����(��I��i�V"O:�x�#Ɠ?ÖP�Q+Fy���a"O����-�#8(��¾&^��96"O�a� ML;>Z���cʪ%B�$�"OФ*��Ő�s#,�]��Ȣ"OB�)�K�>EP�Q1r�ϊHMD`{2"O.��Cf^ 
Q�eO�
D���d"O�\Z�� -6�@z���\�D�"O�DK!D��~آ�	�/3���G"O$C���(��d1@a�.��(�"OZ�J`��~Xa�BU4>$RX�"Ojvm6�T$[����q�`��"O�)rE�إPo�0�Y 0"O�����	�(ܳ$��4ߌА�"O
� ��7Ċc���8���Xa"O�P��O7]Ƶ��)� ��R�"O�8��fZ�����ݜ3�*;q"O¡9b��dUq�얋���#"O\p4b�^h��Ĭ�%�J@C�"O�0�F�Y[*��`�]\>Č��"O�Q����'� !�Y @-:m[�*O�bV�S:���߁	���+�'���%���.҉;��H?KF��p
�'�2�B��[ A�R�rcƦy,���'b��S��!�$m(��J��m��'��P�k�2d|�daA��h�Q�'�j<�7��#�h��&`�x���'�f�A��T/��Ueѧ	�*
�'H
��@N�3�0�`�o�q���
�'g�)��j��Uq6���e���a%%*D�����	UO�:UeA�]���c#D� ��+�vlQ��T-Jք��j.D�$��(V�n!��I���0m|*�K�%8D�d��A��>��`L�I
��6D��p�iԨ.� 3*�����x 	4D�����
��A@l�/U>ܥ"b�2D�H��=^�,ݻ����S��A�3�2D�� 0,���mJ�U��!3n�h��"O|�7i֊.@����L@]*�"O6�����F	��ʥ�=e�=Y1"OٳF��/M.����f��m�����"Oeit�\�4��]��E]78��	h"O�Q#�]>T��5�V�˸c�y5"OJl!䭔�M�ё�J8���q@"OD�RW�V>G	�R��!�u;"Ox��+B!F�Lrv�ۻ���S"Oڽ��I�r������}�`j"O<� $�
�!8���韗4N^�*$"OnH+�Y�M̱Qb]�jBJ	�"O����mB%%g��aAb��8((�"O���d!G�5� �E�iё"O�H��J�( �4���	�D�'"OT��b ��Pk"N!L:\�"O���&�Z1��3��̆K:��҄"O���n��L>��b�g�X1)1"O�q�bA	..��FH�jG��)�"O&��+[�$�^�CC��$t��"O�}��ES*�@�ya�X��mт"O>	�B��w�p:J��E�13"O���\9M��y��N�&�`9�"ORm��k�UHH"B�9��2g"Oެ��KX��"Dʢ��:�2MK�"O���E肥d�d@��)�k��y�"O��c$H8W�Lٴ�C�Fv�%c�"O�����p�Jh�p�ŭvl�u�f"Ot��V ^<-4�y0D��{e�I��"O�8�DB]/Z�V=�b@ħa*�	�"O����%��Q��yA�{Ű@��FP�< 
ʒ35�x���3/������I�<�GɄ%�i#"K��L8���IC�<Aׂ\B4Sq��8�
�F�B�<A�O;+j��1���s���~�<��>	����aD܄]~P�!L�z�<��H�;����i��n"�&N�p�<yq�υfs��4 K���v�<���+�t�*�
D2Y�q{UE�r�<.Ml�A�5/v�gc�d�<)��}?�4s��[Uh�{�e�G�<���8�j�;㋎p�-�`K]�<��f�3Llܹ�l�U�R�<�'�R��ј�&Y�N5L��J�<qŁ\:}�B��e S�Z#�P��*I�<� ���a9x0�6ǘ�r��@�RO�<i��Èa�2T�-Ә7{IВ`KO�<��J�F� �	��ϛ/	����%	p�<��D��>Q�DL�86�p醬�n�<	t�W1�
ms�F�N"4���G]m�<a4�W"���A4��?�jpC�hk�'D�?�OXV��y�aY�Dt��U�?ړ�0<�`��o<d��I3Ni���*]ѦqlZQ������'T�#�H���D�5�T1�yb��2�j���8��8j�E���~,=�O`�h'A�p��ìW���LI��'0�'�>)z�!S�<H@8�� J9d�
�'(�0�P6ɸ��eд:�s��)�S�4lú|��%@S.S�%��<d��0�y���iB�}KR*G	*B�"sFE���	oX�̑	��C�>0�G.�?D��;}��'��	'N���]+�&$�A�I<^(�">���ĸ~2G�І5� �2S.���auk~�<�cnR�P((qGݶ.:�x�Z�<����3� zL���M�q� �i��ɏ�
��W"OQ�l�4#�`Y�S2[��:�"O����H�R#d�����[��'��S�\��)�A	ֹ�ܑY�k�?���
O5yef��{`�9����?.պиf�'KqO�`�W@Q:I���dŎmT"O���1��;�dan�h��E�7��cX��³!:��	2��(?0�\r��&D��*�4���l�1	L�)�eE�t�Ī����	�|�R�{����1�b�bLX-|.��d3?���X8
���{si�Ch4�$�N�D�<�s�'w�(�*��4���%�S�kR��}B�xR��i��i��@ ��S5Z�̒��7D�TRdͣ]n�q(�aS	w����<���/�S�OV��*�ɈWdH1as0{���1�'��X6/�z�^<˲�ūr5�L�{��'\����Qþ}�jc�R�+�{��%\O��p�$�f�zTȇ"�_���5Od7�Y��J%)Z�FJ�x'�͸Yz�C�Ɇ ��xP� �Zw$ q��
)햣?ش�(��m� :C�v!�u��Q�����"O֍�Q&A�p�ؑ�ʆcz��"�"O�d�ui�6�b�1�:/z�Xb7"OȠ�R��
优sҽ�|��`"O>\��i�*/̬"ã� ������>��f������75e�Q�MX"�\0�ȓ#�F���L�<;i�!������ȓBS>�3׏�5�D��q�[��lD}��QZ�y;"e/
�@�6�		<C��%,�(86
V0""�h�6�Pr��C�	�Ë́�Bu�.Ed����O�~CfB��B���k�<T��@HgC	���M��$��-#U�!i�<���Ă
�P �ȓ^��D�c��0K��h��\�.E6��#��:�#�%;�xh��9��݄ȓfu!��]�B��Dd�7Sផ�ȓ+O�u��>Oql��欏Ez�(�'�	^��h��t���"�K�k<�a�F@�<1��C�Z9�H'��,hT�5a�E�<���Y8U�~�Q��M���ո0b����'z��l8tf�
^`D�SS�@�9�`  �H>D�Xw���j���� 8�x@�f>D��ٱ�T�+^�	�$� �j�U�@/D�h��M1d&�8��oްq^��qE�.D�X�֤�'k�2�JC�;��3��*D��rTEP�p�l·!^�B�i�7�<D��Х�P�<�*��I��!ڷxӲ�=E��4�*�#"	�'�!���?7�}��`z9�%�F>��p�E�A�Q�ȓ,�� �F��(� �@$O�Fd�Dz2�Ir�$�Qa)N�rB��>GY���0�$�y�鞱&f]��b�+O�����L��y�jX���	�ԭ9>b�{����yr��5]�.�"7�3������ރ��D#�S�O`���떠,����R�@6���'�9�͕e�~T�צٓ7i|xH�OB�D#|O�y!r��z��9R��}�����'�	�;�F�K��^C���G����D{��9Oh��"hZ�;j�2��Ё7G� 	�"OD���EzD<Cvk�FK���6"O��˶M �_� ��R���>ʍ9�"O��� ���_�H�*�ᏗS%Z1�"O�J���w`거#}��X��"O�&3A�H�p��������"O� �Ԃ��^E�I��A�TȊ��4�J������1p �9��&�@?�`$�$D��@C��@p4`�ւQsxU�!D���1M�-r��1B �yNrqr5'�O�C�I�+E^d#uBF a%��;�gU B䉌Fl:ɂ��L�'�H�+�A��ļB䉟H���G�(C�n�ӒB���xC�I+2`��7`O=6�)d�H�pc`C�	�
��4:��&"�&�r�G/M� C��#��0$�:����l�0�C��1u�s�OX|t1�%�+0��#=)��T?����M�Ti� Y2a ���K�<с���t��H�MI�h�Ǣ�I�<�`@*�r��.~d���H�<�5C�'9�d-� 텫{8��#Am�Ʀ�E{���i+fH�0F�%1D�#��H�j� �!�)��<�c�B ����M�z8����K}b�'�Ɯ�U��q[�4�'F�8]��e(	�'�֨��!��ƱRɎ�S�dt2���I�Px�AqΘ�	��qA�"GkG�B�ɜ.���Fa[2�]	�gW[�">���IRj�0a��iO	Aш�b���,D2�)�'t]�y�����<�5�N%_�f����$7�S�����Fa#�R�S��!&����"�O�a���2@�H��"¼�!��{�'��#}�'q�(�����Tӓ)�H�X�k��4�#<�02¨��!HP�֤"δ��V��̲�냨=]������'t��y�'~D�DyJ|J+O�3F�y!��ْo	5B�]��Aj������w;�I�Ղ�&wl�)k��ԝ��Q�	|���D&6�(h���xw��Yŭ��p?q�O,-��V�4'r\{���]�l-�R"Ob��i��^C�� `�S,jy4,�"OR#��FFD���G��0�+&"O$��wjԯJO�i���2 �0���"OvM�M�J�2�3���g5�@{�"O1�&98���P@��9�S����'N�8�5��0����4���o����>a M(`J�y ��pq�Ek#I�FX���O�q�$n��l���B�$��<Hɗ"OT	d`�/t�r5�䤘�C��l�P�Ol�Ę�h�.�+R
˩8�f8q��U7K^���$"OnR�KP� ��%���DQHI0�>��k��z�$D��	Z��_n��ȓF��X��Q�[ᚘ)��ˡ`&P��ȓ:��X��_��t���V�6�L���b�	6z��v�ҧc'�P`��1_�pB�ɫ	�+�bɺ��OK7��B䉃;��S���xWܴ
���2M2��d�<A/O�,�7eʧ�T�aE˒1���D"Op-8��6:N�-1�_7$�����In�O#��{T�ĭ=����KJ=�$��'>!�	���ъ'��@B�a�	�'����Ì���rp�6�@1�i�	�'�*�BLaJ��*���*�>`S�'%fdyۢ:���ZVaޓ':ȍJ�'�DY��&!;����ýod֑��'c%C�I0G��yU�:G�%2�'�M!�D�Ce��!�d҄!%���'�jl9ǭ��'0�E��@D�Mz����'��y���0��L���E/|��	�'��@�c�N6B�Hq�*�&r
���'�,�1� M3��q!T���xr2��'����c�1o	h�����+eq&����� �08e� 3@X+���{���#�"O*1�S�W�JopĢR�>uB��4"O\����_7wV��N�
[_v�[1"OH�H�c�Z!�#7r���C"OB\zCj߹�&5��ͬl���pF"OD\H��[}`�P��(YP�,�ѡ"O ��� �s��J����bU3G"O^�$.N�N3ᷧ@=G��][C"O&t� "�[�<Q� �pO`�c"Ob!��EFv�n��e@Əp,^t�Q"OұJ�"ϻ=�r�9��_�B+�0��"O�9!V&k|�������L�a"O�u�1��X�������|�S"O���QCB�d�:	�c�5vx�M��"O�8���@7!pd V�osB��"O������isBaa.��s��]� "Oƈ{C5}�.ԙelЧH���X&"O�D@��P�W�B�z%�ŕz���Jv"O^��խ]< ,�ĲB"��p���'�@�c[��і�.yZƥ��y�����1����+z�ܱ���Z��y�h� �r�acL�w��`�$�yB"�n*�P���.�-k�B�$��'!�C��'+��hFS�bƦ�Éy2��	st
������������y�˓<7���Td�  3^�x"�ɕ�y�y�Au�=x�0Fh���y�lۮ\�4���Ϸ�Z�F�@�yB*8Ծ��5D��r��\['�Q�yB�͑e�e�fj�-uȐ�'�y�"ẁ�r1�+Z�|�u��yB�P0	��ڥ`8`���D���y�/�����p�R�Dd���y��m�ք�u���gD��y2#�V���+֔<o���f��	�yb��P���g��|�>�ٕ��/�yRCY�
N�ѐ�JzT4�uo�y��IĄ��jM���Q5�yr�S,P R�Q�T  �<��T���y�-�	+��0e$���`k��yBc���!�#�
��T�����yr��5e����
�UD�h3�cե�y�)O%{�܀Kt��S�@)bb���yF�f�H���#P�Ti���A#N��y���W[@ !�@�x�z�{B��y�+B�K5J0� Ɓ9d�Thzr�O��y"\ h�@p%�O}h8qQ�Z�y�g�$)�NE�C�����,��y�	՚.��!�E�Urp����D��*���"}ڢ@VIT��ajޥ�hxg�n�<�C�Z�q��L"}�pmA���i��ٟG�v��
�H>LH�#�g�r�	E) (S$-��	�J�n� !�!'6��if.�(\t�����`�!��M�/At}*���Q1<]�aHJ�5�Q��¢�%�>yqgO��8\�����cMʴWk*D��x"ʒ�p?���y����������A�ї%qO�>��S2�J�S��!e8����)D��1B�K���T�$`�Qɱ��Z���'K����Y��� Ң��xQ �)נ��4�O�rq�E�`tX�#��|�648Q���&�م�"�rD�D��X�V0Rѡ[�{�\��G�Hh�GəN��)�ЋC�b��q�P��2I�I*�P�4�C-��C��/=��,�#.�6%��`	b@��C�	�;���5�17�Ң.S�<p�B�)�   `�fۢ
�Ї�؏G�E��"O���,S1��dE,_�����"O��+�!��j$J���˖�ü���"O�P*A��j��u�I�R-���1"O�u�u(�B<;���>�6�;s"O�PQ���LRRQ���?C���S"O�jg
��i��%���ѲE�YB "O����.U2b2j-(��G"dm:�K�"Oe�H8t~��v�9oF4�B"O�d�F�ϴ!u��9WS>4R��9U"O���A+Ʈf���Z��zE��"O}�5MF�RL�� ��A\eٕ"O���DJ��99!D��G� $�T"O�4@�ņ��$�Tdأ6�>��"O�8`�I�uI�4h������:�*O��@��Sj^����R�O�$�z�'�,�gA
�����SB�J�c�'��S�_vl�U�Ǥ4�l���jQ;4S��y)O�8��'7�3}�('�0B0���P2��[���Px���.9��YbM�{� \J�Ċ�8�b(���X$��ԩ7LB%Ia{R������LY%F% � �0<���F0f�"!* ��Z� ��J����c�[�eL�EY�$�,��؆ȓY�^{�jX�y��X9�!��Xo�5�'p�I"Se �JGh�ц�֠U��
W?A2�M�G���R#ئ �K�$"�(S*T>�y�⃺Xu�����'Z�,�"�� D*2����/x��$z�e�.��P�BûZw��Ӣ&X�$��y'�ӱN}���C�L�(���P.�p?)��NM�0��RZ�T��
���`���eI�	-���W&��[@%���2̚$W��:��Đ:J�n��!lS�Lx������1k��Bg�߬5<�u���[8���� w���[��D�>�#F�ʣ�ʌ0ǜ�$�N���kQ2g��$ �'ޔ8�i	�0����-̋\a~U"�'���(�i�"�̜���V'֚$1��	�2������Ymfer��	`�ܤ��A�!�P�QJ�8]0���'���H�KԨa��	B1��B���i@	 �T�*�
!�`��M�����T(a��baHF�A��!�wn��p�ř�v>�Ԓ��\�D����F�����#�)�s[�0�����xd��{��ɓ"z��0gŌ��l��8w� yb�^
vQ��=1�#	�i(���`�]�(���1��x��V�S<���q$~4)P�Ŕ]x�����z2��XbǓ˲���H�⑂G���d����L�z����h�+|T���I���ԛ� H k�4!Cj
�o髴in�]{P�P4z���Y����p�\� U��E
I����JA��M]=P/^����Y�D�$��+�!L��t� ��g��|��e��-
! C隕V��9��
4dV���Q 7��u1u��"h�lC�ԣ,%�W��	¦K6oN-�2aP>40�R�6
-����%X.:���Eb��0�<�8vf��`�����f������-M&z�����Œ&AP\iS*Z*+��T�w�K�^YJ0Qr��7��vEڙK�
u�?�ьȆy"=s�˒ i�V!�dy�l>)G�ᣦ؅�|$ҁ^�L��ѣb�<`�yX����!���5�З׆��f�NY�YGiػXA!�d�A����&7D����^�q(��[1�K�J�M £E�
J�m;'�ʸH����@�'7N��pD_�t/��ׇx:��0pB�9;J�RBB��)���n�}6:�hB���!̋
��`vjB5DҀo�Kļ��c�>d��D"�2�D�L�	���'���!Z+^��a���<�z���
�k�l��\�0H�DJ����{��-[�(��W�ۮ" J����B�H��eC+}��bD;N����	�J� A�ٞ�f��2A��u��I�f~Z���o�t�������Q9F�2'�)�` �K�?i*�*sN�(YPS�	P:�%�ƭ��0�d���6q���O`�:�sŬ�=o�x�b۴bXD�P̑&s��-�m�\g�Ta���
�}z��Y�y�ᐝwV�Z��5��f��+6�h�'pR%#�〿k��-J��2<1�Cj�'5�6z�5@$����q���I�Gg��рi	Vb��	�A�|������ܹ lǷr�B���۹N������,��	L:}���]��h�`�탯
�`��4a�^>ڝz�)��<�=�%/O�q��R&
�u�d�X�j
^�'����pN�S�J��.P-LTU�c�^��	�"ȟ�I�T�"	1�8��Ӌ(����'/�On��$��~'�1¦�W�YjP9���O�+q�?�>�b�*��<1p@ҿ\����[v�a�P?�aw�5c�!�ՃӳD�L�)��-D�\`b��,�<膇��p���U'�r�B�o{�e)7�d�ZIpɟ��".� �ܩ�;>9SH]2q#v�0���z����	?;S���GyT\q�H�a���3àڊ@!��z��5�\�FȊ�1��p�BH*E|��Th���=��E
g���B!O�8��@�/@D�@�G'.<H�XQ�8
�2Ix9���P�r��9 Ѕ���!��)� �	��k(�4p�w�H`��rw�>�v�)+��d�Վ7 �|���m�Z��Ɍ���i՜��E+�'0)��&[�ad!��],o�����KW�L�0*
�uc���F�|��@O�7��{G�l�'Q��w$�5!�$o/ұ��T�m����
�'_���m٣t���� Ã�������m��'�����B���!F�p(Â��>npҁb#|OJQ��Ɓ���D �/���I8�m�a�C�F�D��� �a~�+��x͸�iD�y�nt#Q&��' �`�)_�5cQ?M�v�0D���Tk���� s�8D����ڽ~��` � ]�m\� ,Y�s?���'�(}�s����Wjޠ�eϔ>q�z�ρp�!�$ϻK�~��F��?c�4�aD�`�����in����'�b�B"UQ6zMH��޻k��Kד_��7n�j��I�j�RX!�i!H���K���p7�C䉢+������*��k8Dǔ���@!d� A�F�Ө9�2�e��e�\�f��_KvC�I"74a�f��*���I$2����#iB�'fF�G�,O𠣳�W�)dZ��ѐ*f��br"Oə ���9	R�3a�K�B��J���F8�3 �8�a|�*�yޖ�CG�P�6XS������P�2PC�� �d�R�8Dk� �yb&U0T��\��L�"T���5K�y2�M� :(�"��4\����O��0���>]Heٜwuz}��o��@�nl` �3Ur,YR�'���Dʜ�{WT��nN�kahf���K�Ɲ�7�~��;�F�+O�O��~� _�D�F�
^��0�c�T��p<�S��" l����.?�4j�+r�L�IǬ&K�K��W̓&Ia{�)ь2/,�8�G�8 �x
����vT|�ԈƵ?>?uZ�4�Vm#��_2���RmZ�p
�<��93���!�$L���i���S��e�C��[�M�D�}��OY>"=��L�Ah���	�^h8J�Rp(<aF��-����b� >g�)@1[�*a.��r�Z-)�ӈ���~���ƏP`fe���&������7V���\����J#r���(�6�Ly��߽B1OH�퉺r㬹#���}��� T����'�z��qH
&-)`�G���'�r`�Ů�t���kc6���]�*�O�`P������,�B�ms-����B�y0#���CX�B��%�p�O���'(+TG���q�N
/�6O�:P�W�ʆq��@B,�p �'|�0)OR4  #A�k� ��M���P�RC��M���	� �n�,�"O��Ї��4�n��*'Y)��m�x�
�a�>A;�gy��_�]�z��̠@p��
M3�y���q���Q��L�99�X����d[^"+��� ��8?�]�6�lj�i���=O���g��[`(��W `�r!+7e�%j�����.E�����gSf��4қe�r�+r�E�(�PL�%>��VБ��g��~�?1k�/D����Hv
t)8v�2Oz)j�' %F��O6�8�jO0��kDB\$t5�Lp&hR�f�f(�$�>���0�gy2bY�� �ԡ�	�pX"]��$�p%"8H��	���)�'/rA��ЬA0 ](v�Iy���bW�y'�*TC�E8��t�Q(�!�N�_Y����^P���I������(�)d�Y�eݭ�~R"ʪ3f&]٥@�A���)�\-��?��J�5X��R�i�+r�2�p$�QVR�xB\�6��'?�� ��Jx�S����[�}�EQg
-���ҕf:џ�Æ	��BA����ԋ�N֪p����R�֬P��D�y����am`:VLP�N��Iy�����B�"5#�����)�'/��`���2��FK��ȓ^!��p�bK@������I��52O��dKɿB�аȄo�I�3�	��Qj����	�1h�@B��V��D�����1b%�$�\��MϷ/��-�ЌV� P�)C�	@%O��|�H�R۬�p�+�)��Q��G3�0<�F�ǂ]\�@��q?�I<P��\ R�Če�q����:�HB�I�"�n�9��B?��$ �@��*�������f�Ûֈ"��!�Hɨ�)/%I�s&
��yRd� ���uIC�!�P�
r�)�y
� Z�	�aT2"	� &D=9����"O�8�'ЎXUa��	�ȩ�"O�eQ�`� c�&�&�K�3S�$ "O�dIg��,X��PB2�W���p�"Oi��j�`�����ꌵ�z���"O�Y�"D(��(�&E {��� �"O0m�FŬz(��N�'�r"On�q�NE:@4�!+J�|�\�
�"O���N
%�h���*��W�0��6"O�0���ݼ�"ٙ!GN�6��؊'"O��*!�x���І�j�� "O��JU㇃B{����\;��Xj@"O�I����� "bK�gb��ʤ"O9k�� CH���p�,�H�"O�s��-|����aJ2�Z�1�"O�hA�ċH}.��L�A�ڨ� "O�A1�/ ��a�e�,:�D�"O�l(t�2A�R��%� L��Uaw"Ob}kA�ܿ����ŭ[�"��2"O�AY��������M�?N@X��T"O@�5*/_l��^&=D��`"Otp����j��|3��R�Oj��R"O�XD�@�i����,��~�X�"O��#�a�>�T�! ��a�RX+�"O���H}�	:�hW�}�Ҙ�B"O.8P ^���X���^8��s"O,�XR �A��c�� A��H"OΤA6�,B�\���ʟ>.�&"OƝsӨ�&^�ڂl�8_��0��"O��Q��O�]&8�K�-c����p"O �!FϴO�1aV�E�pRT��"O���ARu0D0�Ʃ_>kM�`"O��U#� �|)b�!�0(EH�:�"OD�"s�І$��g��'K�t8�"O�L�e뜭ތ�d̫<\��"O0p����@x�/�h��"O(�Ѣ�WJ�>]x� �H��BW"O�!Hƈԕ}>9�T�Z`t
r"O��0��.0�	�S�`Q♀�"O�H�Cg͒ >Xr���H���g"Of�P���TF �1���3%BX��"O�l7�սE}�H���.:��|��"Ond;'-0wyve�N�cJ�0�"O�Y��"A�1ξ s��w3��X"O�qІ�F�#���Y���}U"O29��Q./���R `�.x���"OI-�*�>N�JD ��R��!��Ų�T�n�h� �;_4!�I0Z8J�B�N�5�� x!!� �!����bM�"�x	���T-!򄇭JZp�W��,|
25#������p�scN�V�1��(H$Sm���ȓql��oñ6��f	#�� �ȓ#��t;df��p�*���#.*�ȓnx��S�Am\c�HV�c��q�ȓK1D 0 �تl	@��t�4����K#����N3O2P%a�6<~U��~!���D�A�A2�:w�@�S�	�ȓ��5X`�ۤB�V䲡�?S�X,��	*dypq柸�	�Ƅ:/���ȓ�j��u�?A���ʧ �0B�$\�ȓ>l,�#�����D��h�H���R�L�#�0�,M��GWo�����4�X���8@��h*=��S�? d��B��0��B��FB��a�"O4�aeB&��%�T���?�+�"O<�cPF܏68��YpC�'�)Q�"Ov��s��p�Ҵ����	 �Nᢠ"OX�I�lS�U�� a�^і�E"O(���m��b�ڌ��_�$d�Y "O��Z�H��n��Y���\'/f\��f"Oր�&��<G ���%��1X���"O.�0�-�bb� zE7R�}*"Ob<
�	�8]Z�Ƀ�d�j��;w"O��ã�д �� f��P`����"O�قa��S�8t)ŇZ� f�=�"O�Ps��dY�(�F��(RY��"O�|�0���A��0��Ѩ^�B�R�"O�}p�+ݎsh��`"���Dk�"O@�ۢ�w�<��5i�%;2"O��+�a ?�ҡ��F-=��h�"O� J�bóZBtx��A�-ÊTBD"O��sA��:��T��t�XQ�"O\�#��� 7�)�h�B�d)�"O�Y�wj��n-0�k�T�"O��Q��3`����� �
�D�i�"O���ɀ�#K������,`����"O��Ro���%-Vru��"O��hL.ww�!y5"��h0����"O�$Bt�ɢnJ�if���q��p"OzE��#K���4�ʮa�L0A1�'¬�p�"�DK���vD��DJ��(�	.D� �5+S0#�y��MC�C��1#�D8ʓH��e�Ӱ�H�����O�;��bs�ɉ���#a"O\���GP
搜���ޘGT��2�;
z
���I���)��<������4%�"R�x�� �L�<I���t3��"���n�L��0���<Yw�K.WH�ƈ4\Op��v��5.�K�P�B����'��	�����M�u�N�4�bIć*���97�<�y�B }�Ɂs��|װ!�E�tB*<�;�D�34�`�D7��O��2'R
$냥�! �n(� !�(A�!�ğ�B)$��@� �4�ӃN� X���BC� bH����UP`�H@ܓ<x����^�O���s0��5r��OT��� P��'�B���:��#.A4�k%Ȃ4wA8����I����U�8`#�DC��p=95g׉HWr�mPEzus�)L'���M�6(қJ���*I|��'1�D��u�C�,I�AŞ17jQ֬�0!�����`�D�Z6�����"��4�XI��$J��};a�>����M�J�>Qa�G�'L�J�i��	����ې+�^��I�%6T;@�Z�lA�O�(�ԭ�6@N��:��B���\����N�fXsT���ē ��Šƈ(�	�sX�T푘h'xt)�A��xjPʓFg���%���ӧu7MĎ+i(�`��<�Ԋ�"6�%���"�2T�X�<A��ŇU^��g�)U�X���&J�S��rg���@���H��3���	J�K81���(J�V��H �
�y��B/� ==Թ86H"}~��f'Ѻ&�Z�Q�\	e��0>!�n�9��1H~�'gp�Y�bӵz��L���]B�9��*:}��+�?�l�~�� mȬX�(��}��i���9�M���|�F�+_���@)μ9_dl�������d�%:��`��IV���i>��#Sm~��dBN,���/��|j%(�y�jU(=]]��A�!D�m��ɯ`��'E�}��jɮ�Ϙ'�<a��#^�Y�>x2FC�v*�U��'�4���ϲUJ� �n�"S��8����#	#�(�O*�a +	Ǹ��.QX���A:@�1�I�n�y�ȓw9�IîJ�w<�XCp�D���Rǣ$����F��O.��#[]84�5Kù*���BqOb� _98��Y��
��b4��_�����*��>1�	T�t+�=*2�X*��ĸ/6�yRk�<.8�pj�hDx}2�K�v�ܝcZ�0#F�(�y�Ea<�e�F�>vϺTx�ب��wʴ|�iY*zYP"� �)���X��m �I̢�9�"OB5�ņV
V��LB�t	�"�UYkb��O��*��9�3}2�G1������h�cpM��xB�bru��K
?tq�F�-P��mI�V�?�.���	Y�tXdJ���4�� EՕp������ �ꀅՔ����*7�t`r'ϕ"B�4��ؽ/�!����ٳA�B�{�\p����g��'�Xdȱ�T�d��5D�$���v�����U��������y�CP
Q�b���(� +���RT=� �|��R�����]N��҆BI$0�ÅY��d�A<X��O���E��1�:�CkȖ.��<x苙Z�|��'�
-A�	�]U�8�)[Nr�5y�}���dH�;��S+K���c��&��9@/ݴ_�C�	7|`�5P3ҳ/4u��*�7j�i�w&ق7�"�'n�xG�,OF-J��Z�6�F �1HQ#^� �"OD��I�eT��m�C9N�{$��3�,	��Z�i�a|r��s�*�����/Q��\r6 [��p=�T�1��%��*n��1���#W8�L�����$�8t�/D��ZÄP8g���aΐ#lg�� ->�61{�<���$�?�g	ҍ#x�)X���oҚ`���#D�t�e�Y>���aO��vi��0��Y�-�c0}��PZ���$��2�>8sIJ�Qn����܀y!�ę���z5�Q�1�&�۷� �vx�A��͝�Ry
8��'�d@АH�Z���@�,n�bY�J>�� ,o�`�OX�І�G�m�hQ��'D�)Y�A	S�V��4jñg^��
�'���w{/c�BϜ�b���l����I.gV��wY�-�d*Y�J��)TO]$BI\M��'�X�ҫ�X�@���NBVe��)f�.���eMDX��/���u�ID�@�O��}��@����D�
?�^\v����䍶m�.Ĉ�E��*����Ď/�!�D	:I�8�K����`�p���u��,Zš�a��H���)ͽ(q,X2넗2�:D��	�}!��L��a������@(�?k���d�>q��Рy?��>�O(�BF��bd���iN;c��P�
OV5PI�=�&U ï>k$,Y��ªt���s���0?�&E
-��l���39�vm9QN�I8�؊�A��������t��k��!?��zX���!�)]4,|!�ݣM������vH[vhA�P��	,���P.������2������޸H��\p�ٴK�b�艇�ɏj�EZ� .i��`��(�M�\��|�h0O�V����f�1b�����_��������;xf���V�)NB�I;N�����^����a���oT�-�*x�ɡ��a �"�S�]&0!���Y6G�y ��S_�B��w�68�&�N0/+�YK�i�|ߢ� 7*��j���'��]E�,O"����E/#͂���"�q����"O�p���ݰ}�l��b�l$qIUc�8��=�g7.a|BĀ>5 xqFN��s0b0�ao��p=�v��Cd�#��d��y�OS=8��p��Z�w6NP�æ$�8��Iϵh.�1��P��D��bSO�T���>qa�E<��ȑf�%�'OlYp�-R��@:2m<2������a�d��G�Q�!E�^ C��H�b�Āc5��s:B8ԩ2g��'�|�D�,O��b"N�� J|�h $���(V�,�qb�/Cp�C�>E��J.C��!*����r��֬?,���A?��i���f$��~[�l��@��XFEA��>�`��Z5���J|�[w	Ċ9�5O�9�*��Oiz-�#F��9�y�'�'0�%@fʁ��V	 �ِi�t ٕ�'��1�@�1O<*��{J?u@�bW�~�flCҠ�4{E��W@.��\P��A��5����Qˠ�ή-����gÉGv�Թ�"O��%��w�Ԩ�H��Dq]�bS�4J � [��yT�>E��(<w�պ��0�LT�f$f�B�ɻ/��[Ӧ��U���k��/e�,��J��ٷ`[�A&?� �ủ�O	�|Ce�ͫ_aZ�z3<�O�	�,ɷ`@pb��0徘�3�/)ta�a�����?���\�m�Kֵ@K�}���I2�b��D��7��zr�3�� :p�)Ւw����,�Ы�"OP�RB��1.=!:�$׶x��ra�>IT�ɮl���?�Ѓ戛R:�(�I?
��+ �&D�r�Z�]�reJ�.�:9��L�D�0D�����,�0@Zb��t]F%�@�/D�{��"aF�;�a'(�i-D����c�+�Ő�4|;�+D��Q� ��q{g���6Ԃ�(�/,D�p`[�O������;�fp��+D�z�uB���Y�q4"q��'D�|Մ^�X�x��C�h����`9D��j������THq�B�4��Y`Ǯ=D�T���(h��u��'*n�u�8D��WĞ�]͊��P�ޡ`Ǹ�C4%6D�8Bv
[�C�@I�'�#��]� �:D�� �Ճ"~2�sb(/�%��2OA���Ǹ 3\a(�
�q�5���U0�V�ЌHcϚ�-�n��B�1D���I�O �K��v�D�*PJ(D����V)g���	�l�/8����c�%D�|(��0k8<�"!K�>����%#D�\xf.Y����AȻ��X��?D���q*T�ذ�$�JI���S�/D���1D�% �)��[Z,pB�e,D���Ƨ�� [���FM��C	"���-D��v&�TO�hvo�$1��Q�<D��xb�Խ�$�ӡ�F8.�
�s�I8D�d��AM�!@1i�WèM�5�,D��)�BK -��y"O�& +VK!D���A�*8zP�`�C�j��L8��?D���#G�����<1����!�ɿ6�т� �8}j��Y�}D$b�)��6���`�lM�T	*���*D��ӄjG>
���&��1<�ql3D��x A��{��z�Z�4�,��R�&D� �d21�� �$�;SǮ!*�h%D�����؈N�8D�U���EI�#c!���H�	D=0�D�ԠҾ+�Z���MؿJJz����1<�ɷa�(�	�cya��GjE��7��a��3�yB$� ���<�}b��O���NK�_���u�<sP�Z7䑬}��I�y=��)��OR�R'4O������; �% ��C�Djs��\��2+x�Ė>ͧ��\��2�	�P�F��@"�HH�U�Oԉ�1�|�S�'*4p�ҋ({H�T@è�����^�B�K��B���S�>ɔL�.L�ub"G˖�R	� 珵L�F��d���?�KS�\="'^��̜����#��|�Ĺ���3�9��)��O�{ h0�����ж\�X��^Yp�:�O�� �O,�(v��/_�"�h��չUx@$�bƊ���R	fz�����A��(5D5�tR"@�qE2Šm�K��TKD�%v#<E��F",�2A�\��D��&T:�y���O?�8��݂?P�cA(W�lt�9�& $D���%�S�'�8��&�=D�^Ӵ�7D�t
'e� ���!�&]r�QZ�6D��Ʌ	![�6*�L+,=#�t�2��0DKA�S�Oݺ�5�D,zh�.��4yx��čۨQ��dӥ��D2�'��E �ixHL���?i������=oP�D
��?AS�U��}�2 ��<%�>=�񣋽XH�'H�R���ѯ����$ߠ%OJ�R�?�0|�q$O��hrI��2$���^p?iV`�H���0��-��<��W2�~�ㄉ��u�/�S�<���WO��9q��o��ȱ4�OP�<� ���Y�|*S��Q�I�FOT�<9��N�1�����c�;!4��&kCG�<YQ��&w�J��1��Z��}���FL�<!�J
g���oKi��P@MH�<��ѱ0ӆ�"Bh�@Cnɫ�*L�<�'bj��k�g��%��i� �DD�<� �9�eT�5��i��7쎵��"O���2�ՉH�=+ԣ��� =!"O�T['��(K��Н"�Vm��"ObY�Eʀ�'��	4�_r����"O��ua�xctY�JA#H�:q9"O���B�'Y���;GE�(�ʽ�"O0��
��o}b�ڔlفt�du��"O�0K��	�$O�	�Ĳ[�H�7"O�����)@`$�ӌ�n+�S�"Or�X �\b�R�J3j���"O�)�C�D/��Ղ֣ "ؘ]��"O���� җ'� P���!U���s"ON��+_8|�Lq�MJ]���"Op<���_и�H��� A/ΩB�"O�Xs�M��ҥ ��F�m"���"O�Q��*Z	Ҽ�օ�\&((�4"O
<;T �9NT[Fg�����F"Ot�r�O�i��q ��f���
U"Ofic���o.�}��jH�>�谒"O�<p�l�6��}C�ƃ.���"O,����ހw�>A��6մH�%"Oxi:g�_&,r�4��T���$"O�TY���<ȥ*�k�&�U�"O�Q�Qϝ�wi&,��J��nE�"O��xv�<nv����K�i�б�d"O�袵�,vZ��s�V� 6 ѣ"O��`�����2�Bh�}��"O6����>J�U��B%jHY"O|uE�&u�D�W��y��p��"Ot�rR��@�I Nߝ���4"O����P�u�|uI�O��`���"Ox|�@GU�H�nh�P�קI�8q�"Op��V�W�PU��Q�t�bh1�"O�4��c� �>9��똆�&<ڄ"Olp� L<2�h2j��̬IV"O���VB(8�`=�FI�5ި���"O������^�D����?"��aї"O:$�"��i������ ��x��"OLl��S�9.��9b�1����"Ot8e)]?\R�v�ڞ���R"O� y��� wXe��
T���:"O6t҅��fl"r�  �FP��"OL	�`T+0i`��&��:/�b�"OHd{e�32I H҅�1�,2�"OlI��*ݛ.W��27'O� If"O�(�
��[�d�j�%�(l���Ӏ"O�@��
έ_m؈B��E�H�f}	�"O�����q�QDœX���U"O♚�f �M�P��e�L"&�}�r"O�5	��6�2!f��|�l�F"O̩���	I�����T�x��p�w"O�`q����5}\p@����)�5h�"O,mX��	9|�Q��=l.uh"Oha���'�<��IR,���y�"O<��� �DSb@h�'�y�N�P�"Otk����I�>r�g�6'u݀"O
ɨ7�ŶK��"��maf� �"O�QYF慆B��w�L�V��"O(��cK��@�$��3�Lst���"Ov���%/�5B��4h���"�"OB�y��R: ��İ��܋"O2�J�cK��%����\�|��"O� ��MҬj�r�� ^"S(H��6"O��sn�?7\�����N��"O� �	�@Ók,�4I���U��"O��Ra��L�5+�4���"O�	k#L�V�Y
G,8�0Hj#"O e�A�$v�Y�I��S����a"O�Q�4d�&p�Ab�D�e�B"�"Oܔۓ���AI���G��\]�"O���4�ւz�n�aI��F�䴉"O(l�! �?��Y�r�ֆ4�( B"O�m8���xܪ-����ؙ�"O8���F?4
y�1f��T��<[�"ON\J����*(��rq�D!m�R@�'�'=A��_�P���q�lY���:�'���e�H�-�f�t��H`��'�MĂ׷?5�T��ݤ���'�jP8�'��.�0��D���|\�	�'�0����L� ��G
	�ZA"�'[�y�i ?)#�4��'ٿ !x�K�'��q5�Z�7��[¸x} �'��L�C��CP���&��o���Y
�'C�Q�U-�7M��E��ir�� 	�'�^��\�s�~�����(�'&P|0&K}�٨3#E�[��'���a��rӰ���ўʖ���'wbu��PI�r�ќ
w:���'y>H�E�N݄��t%ɟ��B�'������f�4���՟[g���'}�p�FĮe�2e sAU�O+�	��'���zv��K���02���=��8�'Q�m!�J"��}�f�4?xNe��'- ,���ȡm����§��D�x���'q ���@!8�*	�m�j���'!0i[a�]�tQ2( �?b�̻�'نq;���'ez�ĸ1k�q�'<~Ѡ�ejMq4$��#��u"�'�`Z��w�I�sW1�؃
�'5��#"b�V�^�I��*2��a
�'~��)F ع(	�5� �7��5�ʓ3� �kS��<H�@�j�}IH-�ȓ}���ί�,�Q��W�BI)�����1A���dw`K��ҍcfT��+� �
2n\����N� �ȓ	���F�|�`�z�` z$T�ȓLWvQ �e�9v/P�����bR�]�ȓ~+��1jZ"5]�Y�5�ګv��=��S?��c�OM$��;��)"%���I��<�j<|H����*U�.��ȓ]ڊ��G�D,]�r�3���<L�ȓJ���pW:��Pq�C�3/��ȓ%��iK� 1!\(H	�#2O�!��it�j�@�XO�dJ�E6Q�lȅȓ6:�0B%k�%^>�1����4J��ȓ:�A@���&{ZZy����~B����1��y�m��{��P�B���N���"��Xc�+-�� ��ܨG�n��ȓkF��{&Ǉ�0�2����"B*Y�ȓB�` ff��.�R�rdEG�z�ȓ:�^	!6�#u(pQ�K+��ه�R���K@iB�RH9��?r�ڄ�ȓr\�HI&N�D���jU�O�h��&s� 蒩&%ld�t��A�P��	>N� `僇aB����	$tĄȓB�b��e� ����l'�4�ȓ�&) ���	3��6���x 0��ȓYb0����h�N4���HV�ц�S�? ���E��"t��HшL�J��-І"O:�4N]Y�h����0��*�"O<9�"1CZA�p�>���E"O6��W�M"p��ݳ�Eʚfx�p�"O9 ���*h��Q�aU�?�
|��"O"��e�8l.tT*օ����(@R"O*TS��$-��	���W�9��9�"O�c"��H�8�*+N�*({�"O�Γ�zln�S�c��` ��{�<��`��м@Q��@�%a��y��O�<)�IA0;�ȴ���Ώ:�l�p$"�O�<�b�Ø�\`q��u��ؑ���yJ�7W�)�e��\�0$P2�y�K�H��+ĜA�ZpC��_�y�n�#;����r��;L�< ����y�h�#˖�k����$+�}J�O��y��
ܼ���V�"q�%��Ί	�yRm_8G��З��H0t���f߮�y"JۤEr�,ӳ�ʸPݼ�8@��5�y2bƫlH����	�IB��jWa��y"�F�9��k��%;=v�j�h��y�"��l� 9��.-.R��#߭�y�hˌN*� 	�α{��)�ՌX�y� Q&���!��Cs$b�F��y���"K��c��L�L��jՉ�yR�޽s�N�jà�!A�ص$�:�yrg��y����4��m���y��b�P���+U�-��8��B,�yB�FY�$1���J�J�2�c�ͤ�y���.d���ȳ0�,��r�
��y�Iʉ2�T�y��S@���GN� �ybL%6�dԢ�$���^�
eLJ�y2��
�B$9C�R'u`�E8�E��y�O/%~9k��R� P���+��y��Ms(9𦍎�p�:ԃ4iT�y"O�h�2Y��:oA. Ks�\�ybJ��U!>U*��t��1cӡ�y���D�x§��w7b��'S��y#�-�-���<~/*���. �y�G�	U]t��P�v�f%v��y�Nޫt������D�8��Ҩ���y"�[�Q��{v��x��ԫ���y"�'��%��C�$p4��p���y��d��('#�}��T�I,�y���%6�fT����#z v�����/�y���&���r5-[�n�rx�c"��y�a]-�DPj��]�`H��K֒�yR����t{���0`a��y�I@H?R����sU�)��˂��y��07:4��7l��(t���!�yr2S��0��Ů	aP�2�y坌9���VƟ(�Xɐw��-�y�h���p�@	.$�Ĵ:�#� �y�$߫@c�QlB�SBL��'X�y®L*}&1�V�L�F�M�!��9�yB�+da���bG>:&L��
��y2eN�"�IZ!��4�`���H��y�D�s�����nċy�m2' �:�y��Z�rĝ@ ��V!�'��y��1
���Q��>\$$��b�1�yb��*! @  �P   �
  �  O  �   �)  !3  b9  �?  =F  �L  AT  y[  �a  h  Gn  �t  �z  �  �   `� u�	����Zv)C�'ll\�0Kz+��D:}"a��6��ԫ�7O~�#�<O��S�e�&zC��(����0����'�`�2�#֏(��hK�@C�}Wd���~�Yt��?];��P�?qBTAŁXi��"(��6i����DÑ}�F��iխ(FV���G��nA �b��u7� �OU�4�'X����C�\u�'DtslղtF��`
vi`��˟lY�/	�4����Q�H��M�&�A��?���?y���?��%2ê��"��="D\ �h�4�?���?��:���O��ӯ���O��җC4nh�m��OY.n| ���O���O����<��d؅��Y.@���O�(�i87T�����!�~١�C5ғ�ў�oZ�I<Z�K�+օ�d �3QBv�q�O��W�'�Bhc�?}��+s/��"�L&v��Q'���?I��?���?�)O��D�|��w�r4 P�B�K�zIcS$[�L��0��`F�vmp�XlmZ��MS��gO�F�g�VTm��Ms2l�{��3�Т,���BCEX�^|3��ɩ?�X�|��'c�č!�//,����b�/|�d0�� "}6ʂ��*Pĩ�ڴhě��h�P���?Eb�̘=t�`�
4��9q̪h�T�=�Lh!,vӆ�h��O�������߉]"���ڴ�1��kS��M#c�i�d7m�*�v���\&��H�����жl�	i5��&L��A(ߴq-���D���`&O�@H�)ط�E�es�8�HK�]6�,�`�����64F��m��]����m�\pn��Mc��],\�TpǦDO�h��U�u�a���v N�8��G?��A��T֦���Iťp��$S�6��ân�۟��?��-7+����E�I�������?��b�'����){7�@�+�r�$�nP��2�B�  � �ix̄1��?Q0����?����������R�b�,�'���C���<��wŅ�s�lE�
Ó=+L6�K1,0d�>!%M�!c� ���j@n��ՉVj�#W��O
�$>?y���"��m	��S���!(6N�矐�'�ў�>��&�*��;�!�$C�㵪2�O�t��=tXf���<I8 U�*:��D!�ɡzǄ#|w P�q�U�d�)X&O³y�P���'�t����+�.=2���8r`�h�'���r��>1@j���G�<����'φM��G�X����
hf���'�B�P���%.Rl�q���J_�<���(�$�f�Z�T�j�I0f��MC��?���?q$����?q���?����+`�P8Pj=�h���� �A
_�i2�Q���W�&��2,�,�.-�/���)����D��5�}\4)����C}ܣC�
5i#�<Kԃ��(?֨��'�)�$S.�DHQ@Ĕ4��X#g�H�`4˟v�DuKBְ U�7-�Ayr�[2�?��'���|�n�Kl�1��ǃ!���:�L�t��'���'��>���&[��� m�<L��N�8%��EH��'�v����|�����W�?��1ە�C�sInјc�J.w!剑q60���{��$��/V��6LP�Z�!�d:4H|4a�HF�N ����ųo�!�
Qm��cD7I��A���7!�$+ͪ@¢E�.6�E���Ԥ�ȓ!���Yo�7s�ؠ8�l	�u8V,��Ʌ�p����@�	��|\Y���K��'t�(��џ|��MßD��ڟX�V�L�����<B��4̻%�����@�q�����_�Q���&Nbڅ22���o���)��$(t1���v��|�Ag�w�(���N�'5ڹ��J���&d���dJ4Xp��30�*��Ã5�����O��O<�$+�)2�m@�t@QQ,퐴U�\�B�1�OPunsD���%eϵK�j��"�B�gծ�"�4��'ޛ�dîf�Ol��̚?Ɣ���$KZ(�S S�`C�	�;X,x*	�%��`���/TnC��6Mع����Z��Qc��<C�	�^'�t��E�2B��y��*CtC䉁{��(���7DP�<�$�B�C�9P��X㑃W�To�sQ퀶![D�o۟<��ß�*v�s^(��I���IꟀ��h��b/o,$���A3eb�ߡ:�M��4$�\+�n�)��w�1�&�H㭈f���aq�ԲWì�L�L\̓7+��"6.�D�g̓.�̝����l�H��r	�w^��1��$K%�¡Kw��O4����9q�,�_
�R�%��j�X�H"D����i�(_� D`"�)�&���,�<y��i	6-"�4���i�<����d�FL�SG�|"E�5*��U�����M��?y���?��d���O���~>1�рU'�H"@��khyd�\6*�C���;K �bb��r"����&�A��.��BbV+k��;��Rr�޹��`Y L�����{���RB��F0��c�ߟGTP�A�7D���á�|���[R�C)�@���n4��֦�$�X��'\���	�O"��o�D�ΜB��Xur	Bq��O��d�y��$�OL� s�T,�M�=��#����a� bt�E	R�} �5Ӫ�4�
��և*�`��A4f��AB�"w,ք�M;������J��0U����bJ=N<M�K4k�Op���'�b����f��6X�Af�W�w���h#`+��7�OB�h��:(���Q��Y�>J�q��'����ҷ_}���C�M�(yXD\>RV���Α�����̟�O(f����'m����KC��j犜�v���+�'�"N�L��k�P�1TpE�i�1�ʴ�'����s�@9���H;~�� sF[3N���A���0�n��vڰ��^E�@�k�bp���;t�哬#�8���lE42����7B<�k1�$�O�}ʜ'����0eSŦ�<Wh���E]�<�C�]��|9��G��x�v.��N��>��̅ml0����� C��sC��O^��O��$� `�H��A��O,���O��kޝ!����S�6����I�����/X 2_V�[�J�x
�����\c>�aJ<�1�B6�dݫ�@\:��Q�è�))#��PM�.ZaEYP�9⺐J~"�i��<��{揗&[4t����x��i��'h���~��'�ў��Ʃ[�A�Fq�E��DZ��Ĩ�"O"D�Ab�6X�(b��xԴQ�S[�$���4�.�D�<��h\�,Q�d�:V��\U��"Q1�ȹw���?����?�������?�OaV�`ͯ0�r��pN�B?>�����E`
|r/�2���A�%NN@�"?��fݙll сt��%b�Ь�1-��"5���& �AWF�C�
��)���Q��i����>�I��M��K!8�ܴ*�fPV���ERğL�	O�';��c�^Cv�&Ə)KL��C� D�آ�V>�2�kbkۉ7ހ�!��4������nyB�W"��'�?QUn��B���F�Ј=*����?���֥���?���e%Sx�0�Rc�4n0t#�bS!L(~̓tGR��Iܚ���g��0��,K�B͍X�<�DD�%^�%����":��"�ś�r��t�����m���QB�� ��~���$�q�@ə3p��;�aի���0>�PD��J�� Ð��5o7�Y��`���a�1qH5qU*�a� �x��G�a���Ty�L>7W�'RU>�"�ԟt����`�捠��ںX_���1��ʟp��VF	��+�y�S�UP�$��q՟b�/�$\��݈q�h+u*ƋHK�d�'�4陥,Y ���`3ßm!�4�hs���!���s��� �fY�]�J���a>�����O8�}j�',�	x�*�i��X�1h�9q���'�衙�T�[����K�H[�����[�OsT�`� M7A��pIc�9Ж��$�i���'����=e�hY��'���'i�9�h��cC/�u�$ý5�<YgEZ";D�Dc�	/x�L���,�e91��`&�X#��q_T����m���$(	, 44`x�G�k&�����ת�Lb>�M<	�M�(29P��@cϬ@��2�/�ȟ��'���9���?	��d�$.pQC��=WHq�uԜF�<C��00�b����~�ġ+ҵ�*�)/���ٟ|�'��p�gFD� �^-2�C�.7�]H+O�I�B�'ՀQ���C�]��������:��*D��±� %]��@@�}DH�Y��3D����P�$ 0k@�
E�4y�a'D���r.�Rn�qi�	�;"�P���&D�tq4�и8���.�WOt��a"�O�5��O��q���1 Dӽ#�p�"Oh�	�)[�y.PHcC2h�H�{�"O�,Q2��E��X!�Ͷ,���J�"O�0S#�U��V]�5�ɏ����C"O���C��f��֡��P㞘�F"OX����,u��81 ��<�~����	�)��~j%&K��Ĩ4�ι)D$E�s�}�<���``)BGI�Z�jt�R�<QFm �Y8�3R/_�s�M��x�<�dKޮ=�y��l°��@{�<!��L7:���)����ɤ/�v�<��4> �YJ ��\H���I͟���$�S�O�Ĺ9T�1�ތ�%�S�0X�y�"OV<!,�u@�]�"N�AQ^���"Or�����8�8�f�S�mC2�J�"O6@�s(Q���)b(�:	=�"O��2!J�4���;Tp���nȩ!�D�~��fkT�f�R��ЎG<?��I.�d��d; p���DI���8��m� �!�� 2	��(Ym�t0r'���P� �"O`�s�؉-��k�-1���C"O�I	��]�E���ަ1����"O�����=&�Xr0j�T	,�XC�'��q��'vl�`��d��y%�܀{�$��'(�"䖃w�@k�ڱ�(�'X��b䋾|�V��ˉ=M.�*�'��� ��'v:�Kf�/z��I��'��� ��?K�,��Ǯ�tԈ��
�'�q	0؜�D�K׭��i�z����d�9�Q?�1��R�T����.N���С,D�ԁ5�H����ˋ'I2Ep��+D�8��-�*=���D�TD3d7D�ذF��1
Uv����-$�[po(D��@TD/�[�k�8��1R�E4D��ЮR�`HF) wIP�N��A0��O�h�q�)�JR�ʵ�ܪ'�N	
���<���X�'��5�fK)V��Z����4��8	�'�>��BG,x�r$���&~��J�'&$B���J��
!U>�č�
�'�ܭy�뜹`y�I��HK8��,h
�'|bR������:���$�(�)O�i�'�R"����~�˧�J% �R,C�' |a�q���Z��@��D�ed`�'�fP1���=Nʂ�i��<p��ɚ�'�6XyP�X�)敫$���bp�A��'�� k�
�� l.���Ė[��Q�$�r��h�:��u��a���Q�F'l^���l[���V�L]pE@-��Ƞ�����t뛹O@l�e�O7-:Ѕ�-��{���R���-ζ�`B!D�8*��B�Z��� �AX�{ɂ%��?D��z��� ֞��4��>�`�bD�=�Z��D����;��Ѵ-��UP������y�����	 B��&|�$�B��y"ퟠ.(��D�"����晕�y��Ir�L�ro�� &D��EZ��y¬��r��X�C���$D��O���yB%�����Ȫ1<lQ���?G��a����>�����'W���".� ���b�(#D�4[�c\�|T���ٔHsd��֭#D����K1�l��F)$�4���<D��YUN4V"�*���s2 c�n0D�<��f0��I�&�ð�x��`.D� i�K_!M�TK�K����(�B��<���ZQ8��HT��"h@�K��4��y�?D��I&.�����-V">Y��1�	3D�D�w���!��`� ��y�*\��1D�\��A�sG`=�2)�&�{�<D�PyG��L��<�ޛ1��M�Ĥ:�O�`3�O� 9eeFx+����C#�(��R"Oy��5Ϡ$���ӈ8�8�"Oȥ��KҦ=L�D
P��A��Tâ"O��@E�:#�� т 6e��La�"O�1��©?Pa�aA7���1�"O���\9F��PCC�_�@q�v�	���~���F�Lq`�A03+
�!f�L�<q�D+<� �hU� 0@��s�E�<a3�$W�P�D�rϨ�1�,�g�<��nf�Z����
N?����`�<��W!p xB�H@�
R�s��e�<�b�'aLAq3e�4X0e�@���܀�)+�S�O�"����Mh��c�nePhR�"O4�vN��h�(��QA��nPn�c@"O� 2���I�a����P!ԘxKȴ�"O�1��+�#���{�i�9B�$PF"O>4	پj)��$)Z$O��Y�"ONL��� `m�I���Y'W8=�W�H���5�O�0�����:\��b���i��5��"O�IV��RT:�8S-�4p\݋""O:1��DI#J��5x��X
B�r�p�"Ov(
ǧ�
m�}
�,	h�E�%"O4�y���$pf�����f4�ZD�'��A��'rL�Ic���F�����Ty	���'Zht�Z�LI�'�@t�Q
�'Y��:�G�&�Z��&.�i�8�	���P�ƿ �F$8ޮIw���h#D�\�S�E8+�aC�mO �b�+>D�p�dc�l(��8�ڪ0%ȑ+��=���$G�Dφ� Җ"�=j�hy�]$�y�!��o����[�]�Mq�â�y"�^�I��Ii�K[Ƥ���h��y�֎dN�#I.�hP��y�d�A�V�1�2A���K��K��yr�'Ul�J1-�>�BQ.A�?�2	W����T�`�ܾn�b��`��YC��A$D�$)D��51��1d��R�v�X�-&D�@����YQ%
+E1@�0�#D�l��U0���q����0��5�#D�@�$���Hh]�M��R
=D�4+Bޚ_�xdC�DA�E��̺<f�Fl8�\��M��m� }ᰪT�O�={�H8D����ܨ����FM�E3��ÒYMBC�I�#�z�Fe��jؤ=i6K�2)C��bNk�F2(��-J2�@�uC�L7�݀gc�r.Lp�N<z����ۃc��$֘ n����;:
!ʡ��7�!�$Z%V|����l�%�4���	i!�dǛt3����o�.i�U�t%�'Y!��Q_�Δ`0.U<	��l@V��$3�!��X
��ГI� p����ҹ?�!�deT��B�'FY8 ң�-X�ў�ᵫ&�'�,�t�U"\cxqJ�)P�$`��]�
�3��X3&������(�E��`X9��Ƃw��I��fab|���l��� �a%���iT��?eHj`�ȓW��9�'G�0'�TQ��7b��T�ȓCf�QX�^$)���� ef���::w"<E�D!
(,?F��"�N�с��M\�!��Ɩ%���a'�9S!>-	���p�!�Dܬp���"&�5>�mʒ�^�!�$ū4�p��'I��Dm $GE!q%!�d�E��h�����u���F�6!���
c�pT�	
Nޤ�8@�J*j5削X����D�;��8��])	�bLb% ��'�!�D�v�f-���^�r�!��i!���W���@D���h��r�S�P�!���%v<��g�> >�M��*Z��!���
��-ǧ���b��!��}"�S.�~G�)A��eˣ%�j�X����y��O)@��A #V#HT1(��y҃�=*x�EJ���q+��y��ҿ�x�31�G.PТ�"�M��yL�7X*H�X��S9Wļ��O@��y2*� .px�݀Er@3ԉ���hO�q�G�Ӂ[Xt1,�!Q;(��-1)<B�=8U��pD�Q8ޕ����?h�&B�9S��S��(i�eBt#� �B�)� ڰ"Q�R�$��1RDHS�f�N J�"O0ِ�c��*9���ʎ'�N� �"O)A�Ƃs�<��N�bp�{#�'���ˈ���\��̂ L�q��Q%N�MZ�p�ȓ(g��h0� �;1��a�R%K����ȓubr�@E��y�D��)�W����$�`��� K~R��$��l�F�<��Ɏ�2���aP�\',(�t��<a���yp\��.b�tkA��ey���p>W�:BTu�R��D]	C��l�<���X�yLa�aK^@xtCu Hf�<�"̾60R K�[��;�_�<9��F�&qk`��lY�S֠\Z�<y�&\i��i�/��	���:���Sx��p)��i���hP�����L�z�H%D�Ȑ�Ƭ`b�xqȝ;z�^\!��#D��j�� G+�p��.��L��M,�C��hq���(�'A�l	SaĈ�3}�C��p�;��HSj���Hܭ<QB��K��9���ߧm���y�Aϩ7n�=Ƀ*�[�Oh�hq"�Q:���
/�F@Z
�'�:Ӗ(X(?�& �6���(��,��'�L�dDӳ'�~�@����2���'�L�aF�׿'Ӥ�˒�Z� g0LC�'Ĥ��*��Xݚ����\1w�,��'ݴ��6Eo�&� 鑝x�
�����MFx���Z�s�I�/���D!s ��B䉦C�ب��юBZh}PP��3b�PB�I�yAY��2��e�P6iT@B�)S�H�������PA�$K?-^&B�	�M�p�����0=j��GX�C�ɏ|�C��ԅ��RE0���=��E�s���d�:�"��O{�d:�p=��/̛:� fK�7�q���'�L�3�'���'�Ёp6(��/m�]04͒'����W�ʺ�Fb�R�\H��d2Ha!��u�'����l�6/�)iB�!I� �ukh�	0k��x��e*hC�X��$9��ba��џ4�|JCLg��Q��T�t��(H�)�ly��'�<a���<;�r��o8 � ��剾'���B*
{�
��g��$!W��G�����?���)�J�J�$�O(��D�G�A�9ئꀢhI 䠥��OX�RcS�Z�Ұ���Ll��9ᇫ���d�)Qs�@�0i@�H؛R�� I��˿2��� �J��
����E��ܯ�'>�ѺJ~��+E#x�"C��A7h����X�<i�W៨��_~J~R�Oޥz�/ю5�*X*f��)J����"Od钀LL����c&gާ-���J��D�>!��i>%#� ��#�<��^+���G��ʟ���̟�xG�W�[aX����`��ʟ��_w*��N�Qp�uˀ�K�Iԡ����[S6�1��5��H�c���"w�?=�?��-[���ͻ!�	+~z|�Cp��=�x%R� z�d�S"7�!�Od�O*8�$�����ʕ��)8D��1�΢<Ɇ+��޴�R��<��2U	��a 츳���t���&"Ozs���)Uh���a	{�t���'Ք#=QA�iT�W���LN_������-� �f@�2�4ұ!���ܟ��I��u��'>21�j����H�}�����U��Te�"�قIǨ�V"[U�e�®9<O�
���9K:���`ƏQ]�<�51Y��=���M ]k�LQ6C#<O�1���'Y�i$��H��}���T�z�p���'�ў F|B ٞM;Pu��i]*�`#M���y�HV���$r��2B���e�2��$
���My���XW 맚?y�OPĢS�V�W��k@Iy����D^������?��� O���)1��B���o� l	�h�E�V#�����%�;{*Mj %%� �� ��e�8R0��I�0ycf��q��
�uƊ�j*� P�/�	>�j���|���?9g�Ox��-�:y��GC�r2���dӉ!.ʓ�0?���K�XQ����h�����nLCx��q,Ob��
X��^uk�@�q�d�Q�H�#�Yß���ҟ�O��� �'���0Ia��_d�끀+Q�Yc&]`���=}����
�4�������O]�PPccBU��!�a������'f�4�ח5|H���=<�Q��o�ͭ;4n�O�N}�s�D�Ⱥ�(Ԥ��~1 9 �' H��ğ���'��� l�z'@N#oJ����!.}袐�""O��i2��Jh�s�+��d�G�ɂ�ȟd�q��&)��q���N�R�A����O^���O�ssF܄Y��d�Or�d�O�E���?��ˀ!'�r̩���]�Iq��T�9�И�`j�J�x��F��`���ȟ��X�B�
b
��C�ѳn�ne �M(��b������ �'��'�}�+�%o���,�a�����D����'t��$l>��df�,t�X�gX�(���7�,D�V^�F�JyKRd+W��X�4I��?�S�i>!��|y�L��c���yE�͂&����뀈`t��(�/Z�Rb�'�B�'�T�'�b:�$<�զ�Gk�ĳ�j�S�����_t ĸ&�E4(��84dG� �T8F~�˨]@~��Ċ!W�m��,�'Z�93C�B�j� ���C�>I���pR�wӢ7-�y�k�T�@& �X%��25�e�@��O¢=1���� 2�tͺVdNZ!����.��!2!�D��y��L�ॖ0�
��b�01�I(�M�����E.5J��d�Oh�Do>]���(���� 
ɴACV$@f��O(Y�@)�O��D�O� �J,�<A�r��/u-X��i>!p�eM�| Ia0^}����g&�%�Z8��A<Zb�2ũFF�(ty�'1��Hv�}{wzTi�	ȕ{#�PD|�:�?y���?����dFU���b2H޲$� ���nɟ�?���?Y��?i+����4@bP�C��B�I���S��Tx����4v��v��RTV�ʢM��n�5F��A�	���Yߴ�?������?��'�P�G�q_�$#��R�O ��~�!P�l�$E{"+�VV�@`g'�B1k��C)��'H���x�O�ӄV��s���nX�i�Q钴�
]��4�?��-��y�S!�?��������y��N�]P�Z�u��&$�2~<<y�b�i���5��?O\�P՟�^w�����P��'|F���hT�$��V�	������OB�a�jb�����?������y!�4T�
�椊�*!ꀳ��_'-)�I���?N>�?ٚ'�R��M��|��d��_�B�SB�$H�����M	~n0��T9%��'ވ������?Y���?A�	�Apd��(x����]8=+rG�?���6y�1���y�&J������;������ay، F`��~iXq�i:�d�p��')�5�ϟ���O8�)G^kd�� ���h�;�K��u�Z�Uhf�i�O*�C���yro���ܴ�l�P�E~��I�Θ�>�8d�AG*���?O�-�Cy��l�Y",�ϓ�u'�O��T�+ V6�x��7%-�eǪS��7�J�6�	��\��O��)�OX扦=�L�ӆP���*r��:z失�T�\#C9��o�VJ�����<a�4N��$�i=����~���l���N��w�����nK)(���� "OR�r�n�<aR�őv-�ym���ѼicBX���	�����<�.���K��!>b<�� �iE���O���	����'��a�O�9#1�:3�u�A�[y�b�)�}�|��(	���j+]�ޒ	� .�r��C�I�v���$&�'Q��8��W�`��C��`x�bf�9}k�����/#_�B�I�f������6)浫����:��B�I�|s ,��"���I�ZC�IG]�U`�,V���ܘ�(V"N4�C䉓W� K�ϖ��\$�ӊ�"e C�6ͪ�Y�gJ_���O�3�B䉹g� \���׾O����	��p�bC�~�5z�ŮT�re�z�B�I:�8P�ÆL�H��ӣC]���C�IL�[��.����f>�bc�`yA��1ZFi�T�*�4�j��P�lCu��c��7�w (�ghڔjcB���{�������{�������'; Q��Ch���oՊV�Q�rOA� #�BΨ"����F�)����
7?����k\�`��q�L#H�*�$�1�0��'e�I
{A��8��W8�j���*B xB�	g���z�/�(h�ya�R;4��C��6;|IR��*u���b2RvC�	8&x�+��5#[�|FLC�GOC䉒~���3mƶzx��sA�(C�&C䉂A�T@�V*�(�4�hB�|I�C�N_��q!,A�g�����L�gI�C�(��� ��"DV�i��
(0\�C�ɡI����I�h���Eޑ�C�	><�R��tn��Te���)o]ZB�V��Tj�児����TDFd�\B�ɵ=�,�� ��,���K&l	|!�D�=֔8��Ίr�ٲ��]UV!�� �U�3�Q_ƅp`K��&�f���"O�u:Q� J&��D�3$�@�"O��ct+avd,��c-�73�֍��mh4!p��<䎹p�Fx�έ�ȓ�d廄ȇ�w}��C�F���L��B�t��)8�'+��ȓo�i�J�F�.�X��7�X��ȓX�b`@�ʙ�J�-�1p�%�ȓ2��I�LI��H��,g:��/��D���-�r��k?@~��4#���lbH"�ʲ,�8��%�ȓh�B��'"ɡ@�ճ�nѶq�0��\�2i!��U�%��I;� �y�x���="�hSsa�{���*�;Cd��ȓK�8rJ�y/�M��⅀y8݅ȓ	��(� ��*@!+��l2���"O���ퟮ%�f��R'�K����R"OZ)�/<d�p��7��+�E�"O��Y��
�[U��i+C/��H!5"O��qա��o�޽30j�("�B��"O�ҏN�E�N<�c�?�qz�"O�$�%G@�yO��&H�'�`3�"O.$@�� ;j�B�׎٠O��銥"O2,@ǭИF(ع�m�}��Xy�"O��).u
: ���>���(�"O���LC�gY0aȁɯE�@Es1"O��I�mz�JZ� C=�����"OL�2�k�c���1!L;�Ze�b"O�Qz�f�U3x�G�3]0�!��"O��1um�;b&�b���,9��=�@"O�)�h]�lc��ɰs�̢�"Of��aC��A�r��4�Ҝ�PM�P"OƸ��H�#~�r���K�(h!"O�qZ���)6�H�u�S�jG��ɴ"O���g�$jhA���U�-DT� "OTXh2� ��ak�"$.����"O��Ɇ�&Z��k����g*�i�F"O^́"D�?A�L)vB�^%̱�"O�Ph�#�S6d�(���VX٪�"OFٙ����dG2�e/[�%
T؂�"O\A�$h_�V)#��K�D�ntip"OV�9��^��ȴIȹpk6QQU"O��Q��Y�n��Qi�CLB��D"ONiAƇ[2X�V�a4�	$���ۅ"O�������$��%R;���"O�@uG֔T��5�g� a+�Ѻ%"O��p��H8�� `�#c3� ڱ"OTe�w�T!U�5vGlКaJ��y�kH?�M��HX�_Z��	A��y�hW�Ox����#%bp�g �y��Z9� `3�$F"�8����-�y+�	+�<0�J�	��"�o
�y�nǗwĞ���g�wP��b�CN�y��ʢJ��qeϰszfa�0����y��:p�!b �Gz�,e�7��yR+��V�Z���uBAPw@\��y2�I�G�r 0s�Q(:���W ^��y�`-o�ura���nDI"B��y�@ ���c�H;檔�R��y2�4$H
TP"�[��X8�ȓf����>Z��ԋ��!P�!�ȓT�V��@�C�E����c�#q��Ņȓ,k�D��A:�"�R�Q#g��D��d���qw�Ŝt�*A���)�� ��S�? z���eɽ>� !@�I3�<��"Od͒���|�h���*�1��� �"O��t�*M�h�)�lȵ�:�05"Or�`@��N���ʅ��#(���C#"OV�����U��:0�U�<��G"O�@P��(L����5��z�"O�C����h�aj��/�ر��"OB��m8J���F�=Z�x�"O�]�CBP>ڢ(`r"��S���g"O�E�� �ʼ��@�JԜ��'r�trs��ax y!%�H�$i,���'/�,:4T�>h��E��*�(	�'�Z|��!\<�8-�!����%C�'L|uZ$�d̃���/ZE4\�0+_@�<	#숌L<��'�*
`	"�z�<�IM�I��rc(#����~�<q�_[4�����K��8�(6D~�<y�a �y��23�K�%�b��Dx�<aEe�D)��s��N.J_�  ��s�<�1�I-��|��L
�{:m���y�<Q�m]1vڸ���K��hD��5�]�<�#DH%P�~]
7I��jVB�Qa�]�<��`T�������Q=��Q4��\�<iW���^�J�8�DӹX�f��G(p�<I#��)=d���g끞�5U��R�<�AJ]>��%��'��=YE��/�O�<ID�ň ����u_8��c^G�<���V�)FV�rP��1
E�(h�@�D�<)Í�ks�Q�'��w��Q2�&~�<�E�>&��5�G�ܧ]aX�����d�<��N�%3pX@�GVc��+A�Yk�<A�,� K�;�	����I�j�<�Rf�Qn@]�w����h2�Qd�<�e$I�]괵@���>$���K�<�r,�ڼ�c��r>�1�LJI�<I�hЩ{\
���
����ha��B�<y�(��z�8��c�7ղ����@�<�Q˕ZK$���B�pec&��@�<�G��:gi��� �Vt��*�-�T�<y#��w��IC�O�0�H��� y�<	��Jk���֩ǤM	���d͂u�<9�j��}������͠�lR��Mh�<�%M1a��̒�b߅'�.L�u��y�±
"<�$��^m�Pk���y��	���y��M��d�
���y"�":_�xb��MQ��(i� ۜ�yB�7Q�#g""[�^�RE��y���F�v ���Zc���D����y�M_ N!P�K +��t����y��G�CH�&mL�1�(TqIB��y��,*��Ga�"ik@gO��y��C�5�r����`��\� ���y2h�3�qSc�Q��Ha�Gܽ�y�"=^�� ��-Q@��R��.�y��E��|ؒ�jӁ�P�Y3@̈́�y�j�`��蝛�Mk����yr����0�[���-!����
���y"�Q�D�6�h%,I/f�h3Em��y�J_�/'�̛��U���A
��y��vUL�y�HׇN�q���W��y2�BW�ΜK�&J�Uy\	�F�� �ybcϚ�p�M�H_�43���yb-V��P	�G�T���C �T��y2�[�*q����R��t�BB��y
� �AR !{4H"����QH�ĩ�"O��C��z`&�"(�;G@�=y%"O^U��Џ"����1k�"1�"O���m]K��`�kR�c�!R"O�A ��B�m��|:�e�#d|��2�"OD�I!*
>(�a##���J��"O���Q!`e�u��L�P*���"O���ìJ���=��Ӥ�r3"Oh��	�X�ViGLP�-�(��"O�S��X>�1 �|��B�"Oh	��!�2Sẇ+r8�!�"OD���T,0�*=��$�zn��"O���t�N�!<Q;t�ܞ[YVh�Q"O5�[�N�P�+��pS�,�#"Ox�9���#M�d�WiM�n���"O|��ALJ!r���BE�@�f"O��hWɒ�c��*�H�$�ԭˡ"Ol�����f���h�5}ɼ�c�"Of�Iϲ,�����Q�h���y�"O:!�����^j�p�߰�x��"O��$���~����SiS�q��*O���I$l֚��`� S�����'{̈ᶪS�V�D|he�۳_�����'�d��c��;.g<��oY���!�'M*��O?Z�� HB�V!��	�'GvqX��QwԆQ�S�ZE�}`�'y��H����KZ�1Ч��j�D�`�'�H�$�-#�Ĩ�f؆h�t��'� �+��
?:�(�2��c^����'��@p$)������cϞd:�'n�%�pGnV�$�a�ֈ`�z���'~\Q�p�MO,����ث����'^�4i��J&/������C\�C�	�0u.��͕^4�lz�(;Qd�C�/2��h0P��=��(��T'�C䉎S�P�s@����X�_"�C䉵<s��@�*�� r��cT�HepC��!#�H�{�A�R��Sc�#\C䉈7���¤�;4�N[ǃ�0xRC�I�:��-��+�>�ib��>�C�	t=H#�1a�Č���� y�C��{S��Y��I�b�|)tm��v�hC䉈,��B����/Ԗ����	�(�0C�I�V�*�����h��ЫiF�|��B��&[�0 �-I�)���r��Ƹ[�C�	�px�l��,^��F��B)���B�I�4���c�P�p���*C;uАB�]=��#���l�@�*pTB�I�u�|jg�l��C������B�I�@��a4��c�\� "ȼB� k���h�~2�TK�ڤq�FC��81�� e$S$����� C�ɪJ��+3&D� T����
@�,B�I/x2d�6��1� Mç�U�U�C�	:�Pi�1&ԕ_�4�B�T-'��C�/}��0� ��7�N����P���B�I�T�H��D}!fhh�- �㞴@�� bJ��C&Ȑ]dR�
3GK+�� 2�T:y�GSZ�s��m'ȀR�ˑ�
|&C䉹. xJ��0p*�h����Q�����d^�'#ZF�,O
 �c�r�$P��o�/@t�*�"Oΐ3�M��|xRt{@���p���W�#X��Ƀ/U�G�a|BdU��(0�u'�oc&9���ڷ�p=���˸	��i���O�ћ0�R�V�b��ާE|huA�"O�I��O˛G��K�JO*p_�5p��$�ot9jD�L�π �)�I
H��4�3��WOFmq�"O���N��rH��f�5a�1�Ta�8n��5'�0�P�<y�EF5�*9����%I)2��	`�<��Է[[X��v"KH�e��疖\�N|����+�a}��iv��EM���0�A��p=Q�l�{�:�j50�ʣD�M��!�boP ~@�� ���� ��+���[U�=(�f��=���4�����ݖOt��gj�=�䡢3OQ�%c!�&➕S��-GވiA�m3>�*a�?a��(�gy*U�@�\i��cPY��N8�y�cƧ
o�,�uo��b�V8��I�%<f}��'h��굊�='
��8���1E��t��'7|��Nҷ`����7��|'��X�' R9R��5�t���C[�l�Dm+�'�rق�˹9�����8���3	�'���:ĪVI>��C�i	9.J��3	�'_�!3P��%d� *�G�)vα@�'����h,Ѻ��c���@�'^4��K��]0�#S��=S�u9�'��%�Q�5��A3$�7��y��'�l���Z����!T�~����'M�e���_�p1J�*�	�~����'q|[R���\��{4d
w��h�'M�,���ɔ0�r����]cx��'�r!c3m�?�
Pƪ:��D��'׾Y�
S @�-6�2�.�(�'�2U �V�tȄ�W5K���	�'����7V5�ٛC���=��D�	�'L�X�炐t�t<� AG1xk
�',��pDN9�D�⮄�Q�Y��'��(x�,���;��vqZ���'Ȣ�8��#h��-9��Kt
,���'�$lQ�p�l�4��f
C��yBC��&	)�)\�h�ެz󉖨�yRM ��
A[p���r�	�y�a
Nx-���F�PK�t��yR��#��V��D8��Q�y��9)Z훵��J��H:"n��yN"�*M��l�	6X8xy`���yb����D
$ �*��p��%�0�yrg�"��1�.�����e)�yH�-0@�����[T(	a&b�%�y�
�O�hQ��`q�!Pv,ށ�y��J9�0#����ĉ���Ս�yrc�#X�	�5��2�*������y���w�
p��a]K`\��y��!5���bd��8i�T��jE��y�Q�WG�ᑃ@/9b��2���y���6�A@�O'd8�`)�2�y��	\R<�"�ǚs�ȩh�I	�yb��(e�Q���׊9Vƀ
��1�y�BK�vyL��2���7����PG��y"J�z�z��=���#���y���%%4����:8��E	ɫ�y��y!������6���YE�>�y�љD� 0�-�C�[����yb��8P�!ɟ�Ĉ��Ș�y�f��Nj���54�4kw'���yB�� qĉ:VG��1+1�yrA�32%�$p۷�F�y�b��h��q�^]2=�B,�y���0,��UP6�֨%�.�� �<�y�B(D���a[�$�i鱅��y�e[��$٣@�^4��0/��y
�  (j�K�( q!Fi r�X��"O4���� 5:0����/�� d��A"OX���y��ax���+.xag"Oθ�bįK�p�R�I���a�"O��*� �))&�	��hщ-�,A"O<�
ӣ�V�~$2��T+"��Tp�"O��reƶ (LИ��\7@���"O���F�§iN@��W'B��AR"O��H��D�&4� dK�G�~ah%"O؍QR!�+BqD�I�����T"OԊtb�"/��$(ܴ(�V���"Oh�� 
�
��A�R�;��"O��A�cF,l�Z��Ϛ.+��"Oƨ���͇t0HH	"�T�p"O q���\�L�Q@����X���"O�<1"dY5+ɔ��D�*d����"O<JV�Ep��X"�=k�ޭp�"O,0:��`��!e!�=�B"O4M�eh	��ǩ?��P�"O�xCR�Ьi�p�zF�Ǵ<� �!"O�Q�F�A�Z�����3x ���"Oh�貤=��������Sj���"O��1f���"�����F�nn��u"OV�ZP�גqn\��Hx���"O��E�/_����ooa}C�"OXH*�� �B�9�I�{�\(1"Oh�P��Q�}��0 ���&Hs2�p"O�C$Ɓ�9� �wO'WF���"OD �d�Ϗ�V��͒pZ��[�"O�$CV�G�F��e�`�'&$~��b"O�����
��,9��M�+A��)�P"O�T���,j�����]={�
�6"O�� ����'�6�XCC!>�L-�"O����3 p������M�0|�"Ob�{�/q�a��%�9LՐ�9�"O`�$�Y�N�
�CP&b����*Oܹw��K�R�Q�H�8n��Z�'0�a��V�(���0i�2���J�'��E1w��J�KwÍ*)�Qh�'�j�#���N�$1��F.'��	�'�^�xQ�P�!�8�CC_-]�pTY�'!�|
�N�o�� �.!���&÷p�j��d�0 ~Z�شsx>-�O��K@'�Q��th1��H��s"Oސ�Ǉ��|�,!i6��n�,9�i�x�ғ˓5dM��ŉՐ�� ��d>hyP �b앯j(��j��Z85raz��_%4��q%�:y3�@����7	�U�F�(V�0����c-NLp��5�O��AU�ڳ0����-�.Hn�y��$�>h.Ty� �Y>�<�m��N|*������[�CP5}O�mq�+�L�<9w����|S�)��{n4�J�@ڰSA)4��e���N��I��)AS}�	�e�ڇ�����\0d͇ȓ$0�
���	52����h�6?�ma��8�N=�a��yi�"?�Ã.QX���R���Z�f�{��@(r��/?J,{7�M�X�t8��:[|:qCa�U, s�0�Ł�#h;��t��;Va�GZx���,?�f��<���5f�As�͑#���y0���x��O���[r��9a�f�2��N�X��A�'�|�i���2ZDD
���1P�J(J2�W���x#�MT� >�Q�����*��'��)
�W�����[�H�F�8	�'8-7�R�S��t��
ެ��T�˲Q#(:��\O�^q���
;U�#?�A.��%���%z=zU�ţAg���I���>=*��ը�-2yDuK�Hɯy�B�IM�R �@�\�T��x�F`�-j3�ԟ��5��EZ�"����<��AR��n�c .΂v�J��eH3I؉O+���Y5^�L���~7h�z
�'��@5���~W�=`��Ӣ{j�}
c�FC��s�#F�8,��JƷ��T��'���� �X8+���P��t:�T�	��� J�����3r0����~�[����<��)�!SK�]#��W�)ʱE~�	�1}�d�עV�"�~�S���0=iS�W�f�
�+�
[����BI��,vm�whא5:�����l����'0�B����B���U��\�H�(�yR��|���) �Th�)0��U��|hF�h4�"@�۟�88z�"O|��� _�e>�{�`�1�ҍ����H��Y�kY�G�V�'�it�"|J5R�H��ư.�p��E�,y[��)D�\���8�^Q����.��2�,m�T�� c�JTR�+ς&���@�	� $�e�1�C�c�p
��Av�\��$�!hK���(.H"��ٲ!epy��>V��IQ�ߓ>�,P�W؟S�D�~X������SX
1O����[��(R&G�B�@Sл�ħ!�L%b��Ͳ;PН�f��ohԅȓR��E�ӻDH�\2�� �n,�B%�T8�I������mڝ����'i갫V'"{6���!�,=���	�'�&��7H[N��P�]11�� �4r��i*��#"���)�$N�4 |ME~����;�PY+��̛idČcӥ\��y"m��m���AK
�pD��2�y�ꛞ3T���̓�3�����B��y��Q!����ʐ�fJ��aI܇�yr�!>	�8 �M���z��V��y���G�qS�*E�r�T�@.@��yf��TP�t�Ԣ��s��;�y2嘸L��!a��� ~(Z`�Ƃ�yr	@�W{n(�&�Z�0���J͇�yR���J��4��g�,N,\x��>�yG,�+f�܋K4�	D��y�@��}״�	iT�pB�i�#��y��=�Z	��
M�tA���v��.�y�)L!�nLJPg��j؃I�y� \�MQ@�ؖ��
��Dz� ?�y��ʫc�ԁ�bn�u�m��
��y2�,3�6dS���jߜ����Z��yB��9b�Uq���4$>0zw���y�#4m�j��g4��b�b	��y�O$e�(�-�[=(X�f�	�y"��)d� 0�`��$����"�O��yb��cE�)��m� *T��j�4�y��qg�dL�S2���@��yr�ת]���Q �w#�pQS�V"�y�V:NG��+���)�l�A��[��y�@S�N��I8�.s����dgK��y����`U�J�"u]����y�;�p)8f�'7���.�yC_�k�����`Gk���6����yB,��ܰ��S�u1�������y"�ǐ ˜�QV�ȑj���g-��yr��2�v�AF@�pDĩ����y򦃷>KbYV�o[�y�P���yrhƙY��6�� #��J&�!�Č
ψMRBmJ&\wj�uCH�Y8!���n� �����<cet!!��(L4!�[�Qp\<���ܥ%�L����_&!򄅝����A&N9*���;G�O�!�]�~�ļ�IDf����T�K� C!��=j����BI�*�$�H��`!3"O��A�O��i`<=S�
�?B<<��"O��ƆGLÆp�gR�_6MK�"O�I1�kϣj�^I�� �-v� "O1r"*�?_>�ِ�P�?��`�"O�1�!�5ʬ)��g�	a���"O��""L�'��	���9#{�I1����7B��K �<`JP���'cF�2�����~��A�b�.Ż�'�0J��T�KD��o�b.x��'�6qrcԺu�H�y��G������� 
� C�f\� ��9|�\���"O����ȃ3[~f��G`�x|����"Oh)1��G
	Cf��Ď���d9�"O��ń��&� ,{ �[=� l�T"O* I
�&Dʴ:�S_E y��"O\���K�&PT�g��8"""O��1����}VFX"��R�*f<�W"OQX`�$�1Q)Q�rC
ԃÊ^�y�bS
�(�ۥo�mbԀ[#� ��yr
F҄%1tG�a4�hӯ]��yr�ζ���q*Y�z�������yM��L����7�Źp
DxR�ז�y�	�!0tEr�jH�>�\5� ��yRKņs���#�GH���`B��yrH�Va�;U��B�f������y�O�Y���Y�9��[�	�yBIXѤ@�W
��+g8��bŌ/�y�#
�E�e��jQY:9HR䔬�yDٶ%���yR�
�E
���o۵�ybOԬ,h�q!�8*5�����y��g�����\�bg�<�(C��yr@�5R� +ek��N��ej�B��y2�>D�꙱'	v�఑�ؐ�y��0h���T )lXF�;r=�y�I
u�\�`2 ���}�ѡ�y-�&|�<P��ķ�P��᧌��y�/C�.J�y���¤|Qx��%���y�B�p4*�i1��7|��REӸ�y�O��+ �r����b�= e����y�O���-�A�L�\[����0�y�aʯ^U�I�%DǶ#WP�c����y2͓���z�+M?}N)K���+�y��56 AY�f��RXJ�&؏�y'E�_��0���B5\T�s�AK�y�*�|e6��&g�91�e������yb(֦]�R쁡����y�����y�i=tt�-�?���m��y���!/*E��)��'��H`�c�'�y"��C_$��Š��u���)��G>�y�!��j��Y�-9k�y0���yҧī7%b���À�2��u{SMI!�yk�"�d�$HY�}aI;�y��Z$ �U!#̐7��4@R��yk\0t�a���h��ݫ1�ΐ�y�.�Q
U	�nSdHK�`���y��}�,J7��a��FE��y�o�K��D)k��g !�ŃB�y/ɇ|�[\�Ot�A����3�y��ت
��)c�/�J��Hr"֊�yB�B>$�d��4\��b�*2�y��C���V썢$�M�tc˗�y�(;13�@����xS�(�>�y�S3h�:�"���+g�Q��J#�yR H����"p�T�a�Ё�Ɗ�yb,�4mh�[ g� p�+#J3�yrR;8K���cP�&��h�1�y2kڔM&l8PCǖ����X��yRɓ#Tq`��
.�th�����y��C7o�|�Pu���Z�<���U��y�/P+:�Bx����$N������y"��>SE,�T#4"�>h)!KQ��y�	&-ܸ�kfj�yD�0�պ�y�D�,a<$�@o� ���y⦌6d���M�J������y
� v�━P,N���x�k�:,ʖ�	�"O��B��U:0��y��ʅ��
m�"O�xda�d��H��k
���"OƬ�cҐai&q	�IB�h
0��"Of�۵A��	Cʓ;�̀�"O(䈃�Ix	��i �o�僗"O��q�D�!z�L(���1@�Ű��'K�$B�Z�~ ISgN4��5ɒnԫX!�$��*,����
I"$6:��b-߰w=!�dP��$�����8N��^�=3!�IrӞ�X�iU�ݾE吀#Q!�8X+� :�؞R�\�r�H�,�!�Ē(W;�����ڠ3Є��5*A21!��G�>(���7��n�n$��	�S�!�$��g�𽺑�г\E��ِJӕB�!�YQnꦂ֊b��U��A�!��Ӗ�C��]�h];w�[?k�!�D�y.L,���l�d��g��r�!�/*~Е ���I�j��-I�*!��8L(���T-3WHٚ�M�%!���V:�+ 큻�8舧��(n!�$��FA�ؖ��Dx�-�6L�:�!�-%� I�f�)`g��a�JQ��!��%!�@cwI��qML!���ܳ	b!���(��B�����m�B/0LM!�d	E�nI��řP�P9*��P��!�[�W��Ց���6i���`2�ڞOz!�G�,X�#@^�`��x�mM�/!��Z�v&d�0r�W�w��X�J�.('!�$�E(��҄�Qx������I
!��@W8Hhq�D^*3*�a&n���!�D��i�z��Bc���l��X�!�d�8��{��B�]n�	b
],C!�$EY������n�����	�iP!��J�UV"�{�b_�> Zl�ߚa!�vF��J2������9[�!�ɵ)�X���ȍ�w�4QE��/iQ!��#d� ���&M�s��!�`��X�!��35��YK�䆆/ބq�ǂZ�L�!��3V���ti�;���i� $C�!���8AM0�s�ӵi�
c�9h�!�DY�7n���yh�6n��	�"O�@+��-s��t�P�СY�u��"OJ0�&�έ5 $��!�
4�T�7"O`p4O.E��h���� ���"O� `��Q/sb��8wd�4פ HD"Ox����Q���B�O@at�"O�ʤF�
P��C�ɪ)Xn�"�"O I��/R
D���I�
�<WN5
�"Of50��.�tQ
$�.n����"O�m�G M-��Uu��tc*$5"O��"�X�Fl9��M�c���e"O��g�I w��6�A�`&��"Op����ڨ	�NtHc�N�\Dl�"O���✂P1`�a剗f$^`�b"O���cA��Z�` �h�](X�"Of�A�H�Oy>d���Q$I��� $"O��@��X�G�68����I��8" "OxEb� <�2� Ec]�/��F"O^(���/YH�S�I�b!�"O���h�g�4ف7���K%�y⩌�8:���F(�AH\l�D�?�y���D��� Ņ�J�R,x��-�yr�0{	�)�ŉT���n���y
� l�!fΊ��x��̅=M����"OC&HA<	���� :~�[�"O\��tGS�]df�`e(Q�6��$��"O4�a�P�u#��� ������"O|d�aK`���P�ȗ]w
�r�"Op��'g��nZV�0��Si���4"O�lx��Ҥ_ID��.�Q~P�0"O�81���i�ځ)G��:��y"O���bӨ_�.�)�g�Y|�Xjt"O<Uz�k�]�Z[D��6��AQu"Oּ�(ۺ�ŻVI\Y!s	�4{�!�ě�W����Ǧ_�5H�PB�_&{�!���c�*I*���P�r���.�!��6A��+�$Q�"�ȴ��Ρ4�!�D��O4$���1�ڡR��E�,�!�D ��~ir4Ő	of�(�톡:�!���`�w�բrS>��#L�:b!�$A�#y�Hv Y�{;��W�$O[!�W��iE��L~P�@f�SM!�d֊]��%sG# �:{<�3��uC!��&&r��#)X���D#T��W�!򤖂.����bN��IlԩҦ&S�J !�dA���d:u�ۂS��,)�]�e!�ĕ�'�2"BP��~ i���?�!�$�
���2�V�0v��n!�d cġ٤
��I���Ђ�̈!�D	�+>=T��l�z̠d�%|�!�Dp���ǪM�j�F08�+�,C�!�րF��;�I#�hk�ꛝk�!�$�&y]J��T��l����diѯ�!��P�$J�j`jH�A{̨�2�ŜI�!�Z�:�w�7cb���q�W e#!�$�I�D$YVĞ�dX�yH2��%!��܃Th�	A$�Y���	q�U.4!�dQ�8�������O�y3�$b�!��& "�rU�B<&?8IG���!�$P�|�ʴ� �u-|d�RM#�!�dŦ5G���'J�$*B�8�N۔x!���>�ȥ�Q�� ,�5I��.Z!�	4/>D!�M˙;L=��l[0G!�T�������SX,���p:!�D��E��� �M*��<�$s7!�d�5+��,r���j�)"��&!�dP�#�VH;���99J Y�%�!򄟋��L:�f8J0R��M�y�!�DG���m����o#`����v�!�d��v���T�G
��)3%�1J~!�d,˲(sǞ�A�Xi�#�J!��53h!�!	�z���L/[!���b*�i*��ؼk�԰��V.�!�DҸF5�	��	N�&M�uB1�٤}�!��4!n�Mq�K�;Lֈ��B�A�!�d�-R���%GCL})��!7�!�dP�`j�=� їGQ�Q ��Pr�!��&���+���)3F�f��4�!�D��X�f��u�F,�m�sHY�p!�$]9�$�1U !8��NX�!�Z�,�(Bd�������Df_�uZ!�1`	���*�B��)æJ�e�!���+�(�p"��z��qa��[�!�$�:1����X�:�)U$�;R!��˙ �N)�śn����IU�]�!��	�Υɦf�"��cՈN�^'!�C�����0f=t2�Xv'ۢp	!�� �� ����@oo�1#f"O�`4bש�ʰ*���)����r"OD����L�ĉi���,W��m��"O~x��gӊe��h�&U�s�IBR"O]�v�	Vlf1�d�9�����"OU��@��H�H rB�P*8H�"O<����Pv��A`N\^�"O��zWY�\���0�j� "O~\)w�ŵk��lڥ�@�Z�l�	�"O�y.��,�fT��`�9L�}1�"O�i��#uo�<{$�țpx�,8u"O:Q�@ψ<��s-��c%��"OLe+�DS18N��+�//E6q��"O�5��Lޥ_>ip�C.52�u��"O��� )�Z����'U�8�"O��p�oTnqZ�[� �{�"Olyj�A��a *���ML�i��c"Op��$��6Q��Ȁ1�ܰt"��u"O*�B�L�e����*2&p,�#E"O�����O:!"`�
��|��d�"O�Y�Vɇ�Q����ζ!��a�"O�%�7f��
��M�q&K��阔"O��	�C#~��QpO�@�$���"On0ȀCN�^����5EЎ.Ҥ��"OXP��T=�R(�I�`�&��"O����.&�,ZM�9�Z�r�"O�a!��6�xE�C=�Z��"O,����"l��6s
PA"O��BAE!���a�I�"O����"O�,�@�7H��|��� ���0�"O�D�&"�I�! �Vu��c�"O��9e�0� ��nC�*lVի�"O�y����.^fL���E�+c��S"O2��O,-���:��ˬeb ���"O�U��BL�[�Z����m�ZI�"O6�Iee�z�$yjr*��&e��"O�ԣ ��=pj��`t"O��2�a��C�4$���AWmh,��"Oy����+�68��ˇ�#np&"O�D���ݶoJ#�*�Q(�"OH��A\+]�,)0T��$�1+s"O��C�9�$q)A	$.�:Y1!"O��3'�~�"!�ф�4�!"O��;�-%РP��N��9��"O�Ԛ�Kr�ɫqEC9� I� "O��XB�Ζt  �˦VZ�	�""OXs��g	�tC�
�1"OP8�
�4m>l���ǎ<
9@d"O
�H7�\�H�
p���%�mʶ"O6T*� ��S���*R?�B��B"O
Di��O�F�G��S�J�Ж"Oz`���Rdr��c R�F�u�r"OB���.*�,���m�4���"OA�'�f���+$ȝ��4i�"O�xcpǈ� *�I��+����"O�\�"N	�`k���R"�	"Oޡ20�$A���D�`b�"O� �u(�(����-!�:��"O>	Q*���-l���B�"O�ܩ�\?<��`ҵ*H=����"O�0�2��./|��8h�>i��`��"O<�ʐg1_\"%��!^^dX�"O����ꇆ����ሀ+@-{g"O p�pE�!LEȉ3BJ�����6"O� h� "g�"�$D�蓅TJF�IF"O�(��n�s��� b��j�<�q"O.y��e��X���ӑ�*x���"O�,1��B�UP�MAq�_��~u�"Or�C��[�l�>�8����D�E"O�EAń�mj%[B�^:i��5""O|
2e�$�b�&HJ8L�0c"O��7%֯���{�ՍKτ�j�"O*�÷�:D��%K*e����"O~ �PIΣ��۫j4@�V"O�{�@�rڪ�㑊�' Ik@"O��#�Ŝb� ܘd,�-k���"O2��'�F9�� ��B�"O lT��!�n(r4I�v֦�K�"Op)1�A�F��r�� �:|ȃ"OR1�a�"�b�'�!X��"O1�� KZ�9z�療4L4�"O>h����5�
�Ě���`�V"Obr�$���h�pC�0�@ęd"O�hˑ��g�t���ѢX�dQ�%"O�IcU�;�����2kl���"O<���N�*'n)ZAa�PMfz�"OR��1D�)Y�v]�����5Y�"O&���@U�MZ!�*G< �PI�u"Ob�1M�-@$�ȃK�FvX$:�"O�����+8s���+C� ��"Opas���0J���5@:mg�|J�"OZy:�h�0d<���rH�SR][@"O�	���W,|c$�ь�
�"峵"OlxF�@5���
5�E�M�p�p�"Oj�Z����2��X�ԃW�lͺ�"O�}�r��w��A@U� (A�<�A�"O��*�4'��k	|8���"Odx�po҈m��	᳌��X
�x�"O�qs�k9,��l�9W �"O2�dn�:C�<��ɅQ�I"O��rV��b�X�@Ä�V,���2"O:�IDX�K:�0�!U�#�A�w"OF�RV%�2}�H@ò�H,$����"OPTHDꄙv�6и�����p�T"O���b��1�����%��z�"��r"O<D�q�ē>nܐ�D�"b��<�"O����iVnhrգ�C�A�.�X�"O�S�b�l���s�[�0iy0"O��1A��1
��3�Cy ��F"O��:�� CLu�P�YzB�f"O�r��M�OJ�V윕_���"O�ir��M�4E�e�C��|�ұ�@"O�9	����5�P�� �.�c�"O��ѵ�N%,�(�`5�"|;"O pX#�R>+9�e@��K��P�V"O �RF���T��g�ʭad"O�Y�M�%(;��3cC�<y��͛1"O�=ؑ�P=[G�4�V��t�J%��"O ����K,K�@trE
��j��0�"O�8���1��y�h(�J�P�"ObP1���N���hV�\�Pd��"O]�N��H[�T�$b��y"�"O���1���r�q��A�bGlMbR"O��3 ÚWՀ|�"�Ut�� �0"O�M���Cc@�C����@@G"O:����K�Z�j))sj^L�N��"O��׃Ջ(���V�� K�v�K�"O>DB�ϮOFȡ'��\����"O� �8Q� � :�6~�� ��"O�(A�gօ[b�°�g�p�Zd"O��F��pqڱ3C�*w�$[�"O�c�iM��~�BԵcF����"O�@��BŦ;.@T*V��?lI� @A"O�zn�.v����
��C "O�@*p�L�3aP�R���W�5�f"O0�s���X��	0�@�L�08�"ON%0p��|�p�I�IM� =�"O�{�Gp���a�?k��q"O����
�4; Ii�o��|f0�"O�4�Ƅ�KbPtn�"v��m37"O��Y����@�͆-V�:u��"O���&��V|xR�%+:
�w"O ՚5d�S9@|���6z&ɣ5"O 	� �?C��uk�Λ1A��"OXY:��( {��S�U�M	��w"O�͚`ax�c��;R��D"O�@Kvd�7@򍪶M���LY�"O��˧��i�\�s+F�x���e"Oh)��)�-ej�*b
ո5E�ո""O��ҧ�M�| 1�S��(X1�:�"Ojdȇ%��%�
P�W�N�&�P�"O$�Dj��!��!� օ�z�"O��Wd^.U}�(�&�0ju�r"O���ǑT����-FNxb�"O]PV��j��I:f�W�!�F�c�"O��
 �sA¤���1v�f��Q"O��#LO44�� �3��;"O ր�!������@jz�
�"O���.@$|�}�&�OX��K�"Of@SrK	0t:���"ʧe)8�"Ox!��O�.�����!G/�%I�"Oε�r�ރY=��2A��ʊ�N�r�<y�� �T5L8�����RJF,ӗ��G�<Q"���w�`��]nS��4aVC�<�2��(K�P� �)��k ��BdOH�<15���{��Z3iV���C�<i�Ǒ��z��WA�JK���~�<�!� w�(̐w���*,�Õ|�<Qdn�>$(#a,I6��Q��n�<YN
�=�Yy�m�阥�(Y;!���6m��Xq���3+�L��7�0O!�Z>O!8I �H2{`�}(���90!��_��87ɌZ���P�@��!�d�-#�B�
2N�Sb�+5DJ�!�dۭ'��t���V"#?��kE ��b]!�D0g�`Y a�K�*���JT΋�;�!�$STDʡ GGH
u~�Q�J�2�!��P����򣓚bV<���#�	1�!�_	�,1��.E&׎d��d���!��r�x	����d�6��S�!��9d�@�թa�"� ����R�!�DB1T �@B'� 8s>��pNVGw!�d�Y`���D!|Z�`Bq_�^�!�ے���H��@G�8�  �;S�!���3J�,!H��3Ѿ���@S�K�!��^�r,����^G��Hx��D[m!�Ʋאp�5c�,jfxԱ����\!�Ď�Z����vč�.,�`5�6�!�$�h^,ѱ�[yd<j'�F�p�!�ę�iي@� Tf�R��X[z!�d|Ɉ��0!�4,\��bI�!�ԜFf�dc�晞}�.�%b��!�� ,��N=��i��NF&J	&���"O����p��Yr'-�-��+�"O�R1�� ��%��L�54-�Yc�"O�q N��V�b���>z�3�"O(��ۚm���F��p����џpzť\56ӛ6�'�V?�@��71����p\l}ꂯ�sp{���?	�&�T��Cɬ<1��!�f�w;l�#qiu>������w8,��!i�F��q�:ғJ���
ʗ�?u�ř��/w͎����;0��-�dӹwmh8�p*��F������[�'Ҟ}R���?a��iK"R?	cd����e" �$q������?1����'���$
�&h��! ��.N ~|��{b�I��M[��iR���_;$�r\P��(.ny9�K��~�IWj��8qQ�'�"^>m ��韘����q�	˾y��i��-mm>l@S#ݝ�@x�wN@�1�����`��R��Ϧ?1�Oi���dy�*%��3Ăъ�@0�iɲ�Ң�ˠF���s�!O�?h��X6
�\��\c�������N(l�`O7|�l��ߴ>U��	=�M�W�i���s�x]�����3u��z6b�^�����O��<�	˓j��K�$Gp��b���`�Gz�iX�6�+�Ŀ~���ųLK*�`W��0Y�T8A�8l���'t�4���GQ "�'+B�'�D�'�Mk`Ċ�o���#FS:�XF�-2)b�[E��?B�H��E��e��mkp�O�Dxb�C��(��1�q���_�i��x���>�F�[�am����� � ���:�x�������BQ�94)����K��pRĈ���?��c�"�?�r�i\����$����'QI����B�����cѤ<�A�'w2�x�c(�\�gfB�BZ �sv��¦��4����ɯ<QTƇ�H;i�Ə��4
�;0�QKz���L4�?���?1�s�Ji����?���K2�5Y�4}�41r�ņ=T)t�Ȅ�ۣ)kМI�e9�h
v���v�b�G~B@��V��0B�udz4+7o� T��P�I,d�T�X��ʨ�M�l 
�����I����d|�uab����K��@�$� Q��ē�?�������4�i<ё��"��H"�b�X��u��'�2�dךO*Lz�V0W����'^�6����'^09���n�B���O�� �����ܽ��Q���f�Fp��oL5*�B�'`�	,�Ģ�o��'�r�� �\���'A� �ʰ���M6X:��%(��TEz"�=A���Y�$��w,��Ǫ�}bv&��U��Ð�<��X�RW5<]����Ƨ���'��7-�OP�'���`NU�b��VEY��T���'��O��Z�#�r��N�*�Y�-�8ϒ8��I�M;�iܛ֌dU�%I�z/��Y�:���	5{,��;ٴ�?�����IWI��d�O�6-�~5��#���a���(�+�'lb�ő禱�V�T�+�a���M	����n��O{kl�.\��B𭝚�<���J>]��&%�n(`-R�g�>r�1�ܴk��ȠI	�@1�k�L�U���H�!�"�u��'Q�8ٛ�
�6�?�����v"|nZ�@J��n�0S:@)���J�^<�	ן�F{��$��J*�eҕm.%����~�Q��A�43�F�|�X?��2���T��Qk����u{t��W�ѩ���O�����<v 8  �   b   Ĵ���	��Z�Jwiď:F��(3��H��R�
O�ظ2a$?����`��4ug���^
��0���V(%��#��Sg����l��nZ$�?��'��h���nZV~RI�13���S�#0>S�]�1��9a�Z�L<���r�<I�I>��j�����,�\X۳�n%�XRAΦ��ɴ��f��2��'4dA!����JHʓA60E�6L-=�,|�	��jԎ��H�(�V˓d3rk�>/�^q�M>)C��.�FJ�*K�wm�X��BP�|���'�9��;�|R�D4&����'0���T��YC������O|�IC���(O^؂J>�s��kw$�ӎ���{����<Aqg?(#<5L�y+�p�@�1[$Ҙ�+��?����I��P�(�j��]�|ӊY��-[�(��'��Dxb� KܓF�� �"�����_�x�d	o�)��:5�	�\X�UH�-�A){�Q����H�m7�	$����s�����gX4 PH�2Lk�X�!��<)�:S���4�c���E�j zFM��Ц�
C���>���!��.1�r�T�N�,�R�K|c!��ʘ'�|�Dx��\P��6" �3b�CH�0�!��WyX�ɡ4��:��	�A��wg		'.�L�􉂍 r��ěxr��H��J��,�C�Z̧6J6�8 �|�i!�a°v��q�G�"��)`w���6 ��Gl �Or�HDC]?H!�'�(�Y���?$�h``eS�~[t���C}�$K>�,]3q{�P�<���*re�I(`F!]��7��u�@́	�'�\��@ ���1�D�P"Od1���&�ꙁf�[�`���+D"O��l�0��
��(]4aqp"OD�0��<i���a� �p��DB"Ov  ����kۖ4B��ڨy�]�f"OjM:������"@�g9��ks"O<���� o���ɰ䇕 
.�C�"O��R,�=}�b4��c�� Պ�S"O����$c�}����8y�L���"O^���D�3e��pb Cؒ��d�V"O~!I��L**L!��B�
��*�"O�Q��o �v�ms�� �{Q"O.�F�D:�"��ɜZ����"O��+H�\�Bl�#��&t��"OBJ�	�0b��JGӗS?DȖ"O�����O�e�΅�$&R�DP   �
  �  6  �   �)  �2  B9  �?  "F  �L  "T  [[  �a  �g  ,n  mt  �z  �  �   `� u�	����Zv)C�'ll\�0�Kz+�D:}"a��6��ԫ�7O~�#�<O��S�e�)���(@ H�E}���lW�h� IVlϊ��@r`�v��
T��?y0a��?�K���] �q�sd������
��1'��#<���/E2JTR1G�%�u��E�b���'��9h�hʷ�����R�h�4<���0<=������OԸp�<v�8$L��՟��������L	�=@<`��\�`�8�kVş��I7�M��N�3��D�Oj�Y����$�OP��"�vIҼ1��Gk9��rQ��O��Ov���O���OA������?���xI��3�\���y��'�HO<�G{�iv���"�(z� �b���;RS��>1�'�Q�I����Iy�IӃ��-:�e`�cT&D����O��$�O*��<A����)}ޡ�Ɔƃ5ئ�2@	�;BA����O�$lڄ�M��i�7��O� l(�M#G�i*\6M�lzj�� �6�D�1�D١A�P����H�'�F| ��i�h�-���ݒ'�Hr�3�B�;�����Z|-��Ҕg��!lڐ�M������?�l�D MV$b����f��
1�M��D��������2��@b�mu�V�Z��Q2VҘ7��覑��4����ܓ�ݡS%9:f�� 5���k@T��ig�F=l� _q�l��*��Ӂ
Ȃk��ӭ��]ߊeXS��3mf)�
;�����X�5*��1�4Q�F�n���Z�,��X�@���K8 @��Yca�L�G���tj���/��L��iX�(ՍK��e���L�¤��'��O��SV�C�a.���F�R�|�>�t��O>�H����l��%�M���?A�EӋe�=�@\�D#���g�"�?���X-*���?�O���m��U�|+'	�w}Ba&1�z���;Y^�WB��0<y��zӔ1���тMK&�_,��`�9��<���ն�DP���<C>��O�����QG�&�B����a�	qy��)��;,sSbHh�:"om���dğ|p�gtW\�zc��}�~��d#�I=p1 #|R�w��q↯$��� /B�A��'?���P�?>i.�14�X�'_��	�'��!YS+׬P/␐��2���A�'�0���L�J� �V�L�J|=�	�'gjm�BB%4`^�)A#"�� 	�'8���
�Ϯ����ؐ$�:��i���'@2�'y�;��'4�'R�w�h����_W�|t�6��'�����p�*9�/K'SH��/��ci�S�?���x���<�F�zQ���6�^X��K_�qK�2i#&�J�ʀhE�����̦.���>#x�`��jx�m2!�^�;q�I��f�6������-O�HW�'��Ԟ?�O��^�@6f-�q�M�jl�'3���O~�d�<��\?)#��?�`q�\�(��E�#��5VZ@ !�O���{}�R���OXb�?�a"^42���I
�$)4ͳ<1���|8�����
�/r)���XH@���?D���w'в$ �2�7Z��+�/3D�|�wo�~���XH�+^I�a�N+D�Hi�-D{+IK�`�O���	�@&D�D��-���%!$G#?آd��"<OfX�eb�O����O$`�1I�!{Ĉ�E`W�c����S��O��Ā*xn���O��d
�0��Z�G�m��s�QY��؀xgJ��t�
z#�k�=O�t� d	�95�H �T`�j��*ƺ&�``H���*[=��P��3լ�?��!�����۴f�v�'�v��g��2z�mgl�r@�ia�'Z��'�"�'��O�1OT � Ϗ�,���,��]��4�V�' �}���xY���*I\{å!���"Ga�!�<�ݴk��ӈ"�O��i Eܭx7"��,M,Qft��"OH���$7��1�U�­L@��"O��#`�[ �s�*W�t�6"O�%��hN��A��SH8p[�"O�=��_;u��ERUO� Y	ƕ��"O�؈�B�g�I+1�[8oS Q��h�X�D�O����'`A&��O��d�O�����VdڃLQ
dk�<:d�
<,��h�Ϳ-��!!%`��Q��d�.M��OE��@�уN@~�Jg�ˬDl�0���ҙ8�Ĺ�7Bk��+7 �9(��c>c�$�'�,F��F#-v��T��o�O��'��%���i	����'�����>�L5�0�K�\�# ��Y�!��	:����о`��cf���I��Mkпi�ɧ���O��I1��E��ȅ�1`3r��"�Z	7N	I�X���������@�]w�R�'��#{�jl�kڃL���a��3u�"�a�O��b��*~��dk�j��zL^5;��7
�!���+~��,c `�\ؤR��+5|bU�!�'�2���Wnz����n����u��4;h!��C�f� ��*��3
�q�͑sL�'��6-<�ݷg+���O� &����`�����s󭔜b5��'b��!a�'�R5�Dx� ��t 3���V;�6-;� �x���7+T@���ڔJ���Kփ%�kw6)��=Xs�Mˑ	Ԕ�M��R���G��[|,Lӳf����(e/�F�O���'����p���=p�$�*��*S�hK�A?��1�OM�w �5S�"�@aǁ�D��)��'3��$��1�.�����sX�P���ԝ\k�\�<8�*Z/��D�O2˧=f�:�l
��S�D�;��
G�\'i������?9�D��I�9#�m��<Q���i�|R� 5_:�)��3H��eI	��d��W\�t�.\/+8���僅��&]�5���S/}m�5Q��	�Z��'eX�S���d��I���8�ݴ�?Y����r�n��h��m�$�Z\"�'���'ў�(�=���$+��b��M'V�v�E�@a��\mZ�4Y�4�?����'qb-+ҭ�)=�	��Ň!(��' ��'�* ��R8J-��'��'VBӍ`]�!��K�{����.�
8�)�'��·�Z\9�T>�<�%@��C^uȮ�	U�G=|��VC�*�\H7�W�D0Z��G ḩr0�D�����d�EI��(����%O�I^�A���O�]o���!i�����|�'�"��_���"qG/Zw�p���-�B��'tfqk��B�t�%���r6: -O�5l�M�9s���'��e�T�8��}:�&I�Gެʱ攺"�\+A�϶vb��'F��'��맹?1�OjF	�&�E�p�D�17��6茈��8;W���d�a��<��+��&�0�Zf��b*�ԛ�@o؟�e͑��:�)�ȏ2�ԕ+ԩ� ���$�O��d�OB��?a��ق�3���=&6I+�"O
�2�H��Sn��2"�%z����|��b�&��<i�ϭl�F�'MR��+4\�˰JC�Aўl�Ү̯bB�'> J��'�"0��,J�ჼD�1Ot|��l��\R&4�l�38R��'�'�N$�1�?���{��}r�Ά�[�T)@d	>�&����w��'9���-E��&�kz$Q�Uc�O�����O\��3�)ʧ^����I��X^�h�� �S� ��I!�?�d�	��@g�	#�&�h���ݟ��'���"�'v��'D�5Hu���n��"� ǳR<~���ˌ�m����	�|�7e�|֌�����$���S�t�?a@��# �`�֤	cT��BN>?A4+���p�'�$;	ؠZ���ɍ:�F�R�Q�H��+�C���"-��d�Ọ}��'�(�8� �"K��	z��ѽ(��PA�'dt� �r8�-���۸a8<S����O��=r��ÏI��m �c��N"!��i��'�2B �]2:*��'��'3b2�<��BEM�Ya�	�|�iۣ#Y��PU�܆#��P(R��-%1�<�%�������M�贃se��%��&iӲ��Dֽg<E�!��+?4�Г��	r�	�P����EQ�m�(��� X��.?Ia`�ǟ��	x�'�:D�'b�F����x�tm�"O�Xu	�:`�,�u�ͯoΎ$SpX�|R��4���0?�Ɵ �RQO֝atvӦ%�ry�����p>12�_�	N�eà����b�B�r�<a�ɏ">��P�"_�{��Kp�h�<!���)	�Q��W&�ֱ2́Z�<� G�	m�%� &ǓQD|]T`P}�<����'ǌ\2v$��AM�6�R8��>��G?y��^� Q@=�EdR�1��h�{�<���5r7�T��Y1&�й��ȆQ�<��g�q���J0_���C�C�<�ԍ��4�6��Pk��;4��y�<ɷ���o�M�pG֓:����cP[�<��iݤl�h�cp�tV�C	PX�'�ؕ�����/v�M���\������$7!��s��X
�l��*A�\�ڬ�	�'�d��F�ͫk-����)�C���
�'9Ĺ��-pЂ�c�S���	�'V��J!��eJf��聙�%ELc�<!v�O�)â��A�y� C�c��5�S�O9d	[a	A=��#Uoq�:��G"O�j��^@P����� �1�"O���@�8E{ #у^|L�Hc"O^�	��		;�5(���ad^Px�"OVu��kF�5d��$���Kp�xD"OnD6b,Yn\�+�j0p�Z�D��A/�OZ	�N�!}}�!���֓Z��"O� ���FH�u���cC@>����"O<)���K5FVh!�H[R�%"O,�2�Ԅs�)����,,�MP�"O�����(�
݊�t�=��'�
���'N>��y���I��J(�����'YVy`��]�7�܀W��b���'8ژ�F#D�Qy���C�'Ed�c�'�n�y�.һ6�^�&�ފ`��
�'N�=�%��-�dѢEM%Ap���'r�xs� ���f��'M6������P<#�Q?����&}:"mBfY�%����B$-D��S'���:��p�Q�SU��5
.D��� O%Z�)j�$�6l$P��+D�L��G�W���2��O)�uK�&D��3�.�H���*��#��![� 7D���b�V.z����&��
x�������O�Y��)�ZQ�5�*�1�|H���2�(mJ
�'��2�U�(W���~��\�'�t�7+;���cG̛G@�[�'�����1��咲��6;�0���'��ǈ�<y�`�/.\��+�'��� KE�)�:QNܨ6�P�-O�YӐ�'$��`��{��A�k@����'��3�(V�,֮��KQ�<�H��'\�tB2�@��>�KED�d]����'�^D��͏�|+tX;���c�"DY�'���p�" �5��\S��6*`��{�ԝ�9%<4J���4a�rU��5)��y������)NεX�F�0Ʉ$��r��#�L���I�AXP"f݆�Ag�cU���� Q�[�)�ȓIxz}(���C���HD$蠆ȓU�`x�	�(yRB����	mxxF{��:���ԉ�pi�,Xz9qA�\�Z��)X�"O�Y�(3����޴bX����"OJY�E�
5�q�%��{N��@"OJ�ٔ�_�=.��(��gD���$"O�ّ�(�/����'�	.���0"O�Ƞ� Q(%��Rl���@0�'��x����Sv�
u0�����6˕OC�)�ȓUS�U�A H��E�Zq�]�ȓ%��x��T�7��P�C	V
S��̈́�U�T|��͑?��mC��� 8�&��ȓXOv���H	6<b��c��(�jM�ȓ}s`TL0!��Pb2DP$v���'?zu`�Z����<���c#L�	�*ц�Ф
�!UOb�a�E��Yt-��8�-�R1��4�IG�@E�ȓO��2�3Q�d�*���E������ ��	6�9r��E�i^|���<�����0	(�K�À�F����}�8C�I�{a�a�ת������Ɣ|�*C�ɐd�mYM�N*Y!3��6�C�	�(#h�s�
 ��:�	� ��J��'����D@�z�F�1Cf��Ɯk�'����'HW{����+z� $����A�Q?YqU��g�R$��	��$�ӄc7D�tGA|a"L�l�����)mx�C��/A�,�A���*��k��R�B��#B��SBn�s3|�B��HrC�I;��IIdl�-58t@�$LH��C��={����P��WD�P��\�2B|�Es��"~��n�I��r������c��Մ�y"�>o/,�ѓ鐛 on�H�C��y
� `�x"��O�Z�H�OΡJ$D��"O��jD�2 �z�΁-EL�ڑ"O
u�C�>і���n��u�D`"O�Mz��M�6Y�M���z634Z�����;�O�ؤ,C2�D B��NU�\�Q"O����K�
.D� �R8��jV"O���D*![�x�a�'��&��h�7"Ox�s���QNl��I��g��]c�"Ox�iWG.	؈p����"�'lz�''zt0W�F�:P�T��HJ؁��'�B�kfB7�Z���I�-b8<r�'^ތY�E�xK��@��Դ
w�9�'��jU�
�ET����߱|*����'�~��r)ş��\3Q(�^��}��'��D�y~6aV�W3�iЎ���y�Q?K��ޢO��X��U��.E�ui.D�Dw��r릜�p �	o�Ȼ&�-D�cVf\%5ƚH��N�}��hq�*D�P%!�-�@<�V��Dvݢ�'D�pӥ�M�!�F�ɗb�qJ��vD'D��$kք
��U %�.w�x|h@�O��S��)�Y��P��G[�I`H���-%��s�'6%[uNMuP��z! "��nfވ��j��&F��6I��z��y�ȓE�B裴�_@ -�s���(x�ɇȓ1˚HY�-��f�`q�%E�6z�І�P�Zm��(C!;B�@�� ����fy�'Q��p>�v��7%�����-�T�p�
J�<�ΐq^�i�וj�(��@N�<��X>-�4�H@H�3V�)�a�L�<�5� ��0�&�7�x��6b"D����UT�����Ҩv�Fe��i=�O��P@�O>�Ek�lV���'�1u��d��"Oj	��nY����F�o��y�"O:(i`�p���1e��Bh|i`6"O�u�J�' Y9���6y��`"O��AGH��]+1��9il�"O&��i�.>��3�]�Jc��@��76Bܣ~�U�Q9,�<�*���( �.�D�<VZ:6o�xG��'FD�!�W}�<�����E<�ݰ�U�����q�<�U�DT�dpv
8Q�8 (t��l�<���E(o[JDQ(�(]1�0*Wn�<	���w7��c!��&�ph�Xr:��d��"~Br@Z�R����tHL�����-�y���<O�lpŋ>F��&�W��y"@����Q���Vo=p�ᐧ�y��&F��|��4dl���H��yB �upY���V*)�
O��y��"D�~���lE�v�HAF����AjB�|"o�<?��g�L$0D.Qf�Ѕ�6��$*&��.��-B�Kӛ�~,��l�0}j5�/{�Fb���$����ȓ,O�\Zt!��f�L�'�*`�d�ȓ�pr�r h�%�'e��m��	�T&�	F��U�Cg^0d��l{w�
B�	?\Ը�D�ʆt��b����C�ɼ8ʹ�'N-�D)#u"��LC�ɘ#t>����V*nHI��TU�C�ɦS[̵�š��7e
( �3}X�C�I�Fi�xa팤 �X�"�Y:�f�=a"D�e�O"��L�q4�;��ʂ-���'�n�9aŲn�����v���)�'�&xB�H��9w<����+?�аK��� ��B��U;/2!'�Mh���q"OT00F�,~.Pq
�
2< �X�g"O�HJ��:��c�^�iLP�A�'�>lR���Ӓm��1p����/���"��
��Ćȓ[�a
�A1U <�д�T8�tt�ȓz�Ph�mX�2h�h���R�W2>�ȓGTB�gČBo<ȴnW��5�ȓ9�Tj�ɕ�
���dMٿ/8�Q�ȓ_g��걍,ac.j�O 9�=�'OzpB��u�gh�GE �3t�R8D�n��j摋��F�YRT�󡛿e���"t(R�h
�)Ɇ�c�C[�q��	��iW�e��
`J؝��_w�����v�~�I�R� �
e�M��ȇ���i2�	7�6��w�G@�ѕ�ͽ8i�C�	$fZ�Ys`�-o ������C�:'��gi.E֢E��.�Qp�C�	%���BC�]�m
W�%��C䉞5��CE�w䖝b�E�R�C�IY
�a�� ���"L�fT��=�!�I}�Om��[c >u����V��&�`�K�'��h�B��2:���Q"�D��'�P�r5A]k��upV�B�G*,]@�'t\eː. <7�ܠk�	�9)�jT��'�h!�S��z)�,r A,Q�\�	�'@�%�ōg5� O�-M�^���.�!Gx��iԅ��#K�sL��+��]6q5�B� J����3y��䬙t�B�I�a�\ �/R���@,�/�jB��"%1ZXJ��N9J��E�҃Լ��C�I�i:M��@ȯ\�ƹA���A��B�I"�81�❒8��M��`٢o�̱�=a��~BD�$NL��'�"�O}V�(3!���H��`���b���8��Q����?y��-����*�����͘��M�2�y�9K���Iʢ�W�0��SQ�'��4a�I��K��B4^�c�q݁��ʇ�["��#iT�e��T�S�&�SVZu������|r�a��27��!���#8�G�ny��'�hd��~���dj2��%�
�fW�	
66�8j�*N�mC�`�U�٨NG��G��Y���?�����)͇n����O��C�I\�X�t"L�8}v����O ��G|�����Xq��$O����jr5��o����0��OS��V�̓B����2M�Oٸ��iA٪�ٕ��L{�c1���1� �`\�	7"���J�A���<#�'9�)��5?a��o��b��B��hĬy�<�E.�%Ik��'ʐ�Vh`��0��u���$�R���t	ET���pժ�\F(r��]!T���'����*�\��'���'���}��I�Kw(�b�R�>W�`�7ʖ`��p×!^�7��IZB#�-I�,U1��j����U7!��g(&J*$	@e��q��X ٤D���/]�� ʖ�,��I0�I�(��Q% �v0fC�3r��'�P ��q̛V�O��O���w�(���V0��8���@T�C�gL q�'AUF���4бd����h�'��6m�OD�=�A8��4�����`ӿt�4 [�g��x`����?����?Q���^���Ot�
.F]� /7T1� ���Q0f$�r�΀{S2�B�gB����L'�T3���1AX����\�B؃c��.LC0�5$ɉ]����	�MCp�d7T��񁭞Pe�JܕR�<��/ړ��OL��V+��� ;�g�dL!@"O@@XҢ  zk�	ɀ��="\عa�X�P�ٴ�?�(O�}H�O�A��OV�S,q�AJJ�G��ss�?CZ�DL0c�����O��$R�8k�Bu�żW�2�p��'t;"��[wǔYA �F6ٸ@SmԲmd6�p���R)a�l���"r=[g�@�/nP���DG�D��_#{3��b�̴Zw�bߴ��O����?щ���qɖ�s5�Rt�HP���$5�O�H�EL�}�dh�� ���s#�'K6ʓr:̈𠮊CMf�P� �gD�q�'u�h���'j`�z��' 哷[����ğ9��,;�q�g�� D��������21-_H�x��B�h\�2�˨��i �S�y�<�6��D��ȅ,K`�	�V�lܚ�	�+Ƕxӗ��N�<\b]w��ΉB�[�TK5N��IU.�;c�3Jq��4�~�'��)�)#?� ���-���Þ*�(!2�"O��1�ɚ��I�B�@�s@xAKs�	�ȟ�������CFQn.r,Zu��O����O쬺�d 2w�6���O ���O~(���?ɇ�%.�I�E�VTM���� }�d�bPh��m����#ܜ�L]�̟��4As�G-
����ؽKڅ��
�g�hs�G%p(Vmz�Fб+�.���'^��,�/��(x����y�z�O��Q��'�"�'��O�S����Qo�0%�S��8p�B�I�`Um��J�8���Ö�Y�;���dY���T�'��ɫ��4�|�
c�B-`pc�¯At|�:PG_��T�	ӟ,��韔�I�|��O��xv(!�b�,Grf���Wx�P`��&���M7a����<y��/�D�jE�ޅ�Ҭ��F`�ɤM\�e4pى�(M���<�M�Ɵ�q X)7.0���xl�0,[ϟ�E{��I�q-�@k2�ИW"<9"� XB��,�Z����O?G���Q��0$�4�A���'�剞w��O"��i>�Kჷ_K��`Μ�z���p�I�OF���O��D�O��
�'��m���<Y����喝k�J-���/WB
�s�'vX��+Y!l�jI��ǱR2����Ͱ�Vg��V@Iꠈ�@�hxE��U�'�j\��wC��%q��$u>��s��p��5DA�sN*�j��OJ��O\�O�@̓0��UAP�(2����݃`{R1��I�M��iQ��Pe �대��Ǎ�4����'��7M�O����O>��?a+�:�:o�lP��6�Č`ai^�����8CHS�{���-e�$$�d���p�����RL|�`o�l�IK��O�$Л�.^�L��nI�;�!#�aӲ�D)��牴$b����ON���O��I{�L�k���<
��@V�H B����ʦ-�	���	�<� �Nnz�̟k�U,H;�,�@ͤ�.��ė7R���?�!m��y����$�O�	�O4�	O�4� ä��H~<@S���N��Eڴ��O��d��T�d{��0�D�?7��6���  ֋eX��y֊�s�����`}�I֟ 0WH���	�O,���~�� 	;+�8b�DB�G��m
�����8e�I"M����O@�����O��	2C�x�s�������l� r�BC*¥+ ""s*�æ	͓YbJ��	韌rPK2����?��� `VUm2H�܌y�(_;zt�A1�Ԟ�yb���?���)��n�O"�	�z���s�rd���U�G����2�F�3��)ӡX�\�n��<Y��^�M��i�V	R4Oם�?��S�W�0DY�ܫP��A,�D� ݴ))|9p�'|&�Q��?1�'�?)�'W��ЙO+4Q��
Ig~���idr(qҷi�^��'��l����I"����)��T�
�R7���]�����Dx��B䉡5n���`�>&T���OQ�f7�O�ʓ�?95[?)�'x哅�]"v�N�Ph��x0�>�Xܴ�?Y���$�<i���D�LX��#	���a���  x�O�O��<��;Eg���s��:+�v ���R�<��GR�"Ӳ��W�ݲ�$�����N�<�@�]1(�NL��--*Q��:#N�<q�o�r��%��֦@E��J��\u�<�1��4$��P��@��A�~="�c�t�<�)��<��PR,K5~X�g\z�<q0�#3%27�ǥ
~��Q�Z`�<1�hi���C��R 1�@Q�!BM`�<�߳"�bɩգ�5&�Q�3#�[�<9�`ٽa�N�d��G#����MY�<	")�I���́7�v5����U�<9��%Xy*lA�x�eBSK��B���"�	t��L)4i����ѫ�VA4:���;e�ġP$��%5�0g'�\��K�b�1�AZ�g?��5�ƨQ���%s|�ٶ�.SOV���O<8a���R��b}���`�&�\q#S�_�%� ���A4f��C���+ y�KMV���>Q�ı"��Šd*kBM!aȄx�<��ECR>�]@0$��K/.tx�ƛs�<�b���W|��Ƈڬc[DY���F�<q��$���˷���>brT��,I�<��e� )�劅
@���V��C�<i�NF0
*<���Z�>6���A�<�lT�Y�z�F�c8�Q#d�<9s˟%�Dp�ң�3�����L]�<aP�Ӣ00.�YT�< ��+�WZ�<A����3�\��`K�%�K���T�<!���S�������6%L �c�N�<٣� `���"���.0`:l����U�<��(�3_.uc`�
�E������[�<� �}�V$�5ԄIA+�Q�>�s�"O��b �Qv��L7P˨��T"O0�rc�$Nհ��R��'hY�b"O*q�S�M u������>d��"O�R��-�*�:2�S�_� 0�"O0 f�h2����
�?>K�h�"O���n��If��!G�u�"OD����+l���E@��-;08�"O�P���(�`����ژ
 ܨ�r"O�!ˑ �9p��0k��$�^�Ӑ"Ox�A��'�����a��F�"O^��"��;� -�� �1&�^D�"O�ɩqhJ�R���K��A3n��ؘ�"Op���
H4B�(�0o���"O$y��<]�<e
�aWTd��"O��Zv(�zW���D����٤"Oz蓫Г ��!N�6{�H��r"O���AΌ@~`���L(K����7"O�p�%��%�1B"̊$7�u�S"O M��I�D�i�C��D��"O4�ۅ��k�Z� �����"O���F%^(ې���±n���"Ox��&� FV��Wl\]����"O<�Bq��&9Q�%Ǎ�J��b"O���"�B�"�&;v$M~�Nu�t"O��ʐ�fq��7m�>c�~��"O�}jD�<�4�
clA�=�L�W"O��qԥT��z�+b	��%�|��"O������.�(!�3�ε!ƭ��"O|��EGW���j�A��	�f�W"O����fJ<4���qD��/V�@ *�"OHUڗ���'9:�������E"Ot1v ���z���M&�Z�Hw"O��`���.Ĉ�Zq�4}{L�82"O>����T4.��͹ �>zA�-�"O*YQs޴{`��k�%2���"O6K��T3�i�p��;
l	�S"O�ɡE�I�p��%۱f%��"O�(r�Ȥh��ek�_4MZ��f"O4�˵���gC`�ɁM+5�0�"O�,�B�C4��#F��3	�"O�ۢ#	1̢$�DF�8���*�"O�Xc3,�,�ĥ���!���"O"�J�&�h�pm�2Bߛ�|X��"O�t�2��bM�Y��NG.@��6"Oa2ce�p&:A*�JŠ:�H��"O�)V$&A�z\���7Zfd��G"OPyjuH�L��)�D�ĵ}��y"Oju��I�C~%J�P����0�"O&����	(|��ЈU�P90����"O�4*�@$,y ̀/{����"OX�Ö�J�!C�����m��YX!"O�h����=n
2,
ʞy�MJ�"OV�*�(�$=����KV�u��"O��1�-��>xn��#�� #) �"O>�k��*w���*��J�A3: W"O��`��8[���F�8,YP�"O��Z`K,/���ۃ��'9�9 �"O��8`�/��
���,_�Q�4"O2|��B�3�$5�g�M����n�<1��Q�8�PzRhR�r�{�*�a�<QDB���9en�K�ܙ[��G�<A�-F6
�{�OCJ�A���MD�<��D���n���nʭEsZ�+s
B�<� ��[�)Y,a2���W+�sl�)�"O����h�-��3HΪfNH�iW"O�H[q��(G��T��h �Ү���"O�99񧘲���e�G���뷦:D�(�r�Y����f�цY�FՑd�"D����$52\�@�
Q�m��,`�.4D���ZxP�(Rr��.l�h��3D������N�=�bn��=u���$�+D��
��+Q�2�j���v �D���.D��b$�
3q��:�i�*J�NxIA/.D�4�2bK+{�`HC� D���#'D�P��"-t6]���ڷ�Tz��#D�����n��	�)v�$��� D�t �%L�;�h}±Nي6��$xQ�3D��U�5[�$l� aI3u��� l'D�H���ؗ]�)P�G�}��"��&D���L��y�%3�CF>CLx��4�6D�@���"�,�J�&��T����!D�K`��?mM��8Ҏ��x��uH��?D��d��3u7�L��Fx�F�y�n?D���,F�RF)b�/�]J@�N8D� ��L�B���s��6kZj�	3&<D���3�;��#�~�����7D�H�4��-\���7��Y�.\��6D���5���5
�a+v��:JO�5K?D��#F�
:'�(l��ڗOw�E��8D�Hc���jW���T�X�V���`!D���3�� ���BX8G�zP�&*D�(S�b�F/ؐ2�mU�?>��")#D�����R�6�!�њ1N�S��?D�Xd'>L��U�&�c4��"�! D���2�X�3$�H�3�ܜY�c=D�X��'^�%�Q�QF:P���I�%!D��Qu�-_��Qs��uVD�3w�#D��{%�*3�QF/W�W+B�1� D���hǣ�����
-@���!D��r.W�w�*����]')�`0G!!D�Zv�[eD6�tꈤh����!D��Xr��4V���BL�,5N���3�+D�|��,�#<=N<���V�H��r%G,D�`�n�..0}��	�,�|�9P#-D�$	���!v��$��Y�T0�ai)D������
�v���D�$m�̨3!2D�0�唉8��)��L�'gZ���/D��F�W�V��3�䜇@��E��-D�pђ�8`5�@�C��yӆ�,D�hz`+��|�ސQS,����< �g+D��JBC�#�^�ځl �|���(D��Ii]4l���� ��EE��ʷ�$D�����%g�8`�d�b��`#D�|���R�EV1P"��:���� ,?D�p�F-dQ�56]���!���(D�d�NHA��+�!:�z;e�$D���R�M��(��"$!p@ŉ@� D����)W�%*D�4I�Dc&I;��$D�����5t[Ґ2�m��O�5��I0D�l���D�;2�����b=�ɇ�2D��@�l��F���[�S{��l(�l#D��4Nٛl�f�#�]%6����D?D�$QF�]�.������3'�\3� 3D�����L35��A	�NS,���@A4D�JG�@�]�U�@��q:j�p��2D�� #Y:/���xA�N�Y>h�TD.D� �@��/U 0I��$2^��9AG*D�� �ဥ �1�
!�`J%Rr��"O�D�Uk��2�j�%@*QT-��"Oִ�#&�=D�:��JȂ`A0A�g"O�Qb� �x^u�T���&Q��:�"O�}����?h���EJMkLD$�S"O��%��/��)Ti��0<��"O�ē�k "P�9G�J
C0���"OFeҀ�4�y�-T�s�"O(�i���X�։�a�Z�T��"O,�k��ˏV>��dN���^]�d*O��� �Ii���fn�ʖ���'8(��$��]@��EM�J�B�:�'*�qR�	K*5}`��tQ C�d��'J��q�R�$�X��"S�@�����'&|��ό3�n���O�/�Z���'����&Gؤk
�B��0fR�`�'k�sp���wvxsR�M�R�2�J�'?�A����y�O�R3�YC�'3��E.�>{,����ǓEp�9�'���<8R]Q� 7�8P	�'�6a2%�Grb$��i"ڝ
�'��Q��L՜V R��C�#�>�p�'����8j�r`��A�~ �'N�Q�A��
�B�N_�wpr ��'��� ��D�u�⡃?B���X�'��y�⚂?&����jZ1�T��'��8�B됼_f�eʵ"V
.pN�a�'�ҙ��S�o����8W���
�'�f���Uo=��s� F�Xp���'w0��CA���#�эT=�a�
�' �ha�W�0X�R�H�Vݚ�P
�'���w�G2iR�}!b�H3��b	�'����`��/]����+�P�Z	�'��8�g�(����óN}�٠�'���Ɗ�mq
q��'O�,�Y�'��-��/��t��=��_7X��s�'�B�#E�j$tx���#@ήٓ�'�p��(	1v4�#D��0�X�"�'������( }Z����S�I����''�����u_ڕ�r�D�~Xe�'Hh�i��I*f�q���	"B��#�' z��L�v�=єjޚ�
�{�'��ҍ�[H���,O:FPv�+�'�Z�Xg�O_�XU[F�./퐡r�'�0��(�6)дBCq�
U�
�'䪤�a�ѡ6�D��R=6o
|�
�'��-��ϖ~w�H��@����y�'.�u !I\�L�V�H�l�0�̔��'Y
I�"�
=C�zĹ���{��k�'�aɃ.�7@���Įq{�|��'����Ѝ��z�T�8Ь��U�a�'q�1`�t͡��Hb��2�'�䚆�Ҵ]��� WH̓ZL,�K�'J�H���9/
�5��$W��z
�'��A�m�;WҐY2`�/O5��	�'0�l���c����ƓL���s	�'@q!�b�B���ˠ�	�C~��P�{��_0�)1�!6kf`W��ˌ2#�8�Sk��5�
Y�"�F�nAS�"�N�<	'���Oa`����'��8;�߳0B����O�$Ο�(��ɩx�Ќ���Q=jb"��A�ت�B�	�5�t1`�T���ܫ��9O���[�B#v�@�x��<�O�H1��t�Ճ���p��
!�'u`���/*B��}�]2�H�j8��d�PC�I�)��Ջ  �w�ڑ��o�K.��۳�کeM��� =C%⋍+|�+�ʟ�+��<�r"O���Ql!Dx{��	*76����H�1~�'��´�<�5�̓HA>1Q�2S�E�T	NG�<���C�	zش���@���d b���Z�>����]�)Ha}R�ر:dԙ*���o:(�cO<�p=)0ʋ�A���j�Nq*Gˁ�a@�#�DQ���NS)�aCF�}�j��&�ulP-�=�v(���i
�P��4�D#Y.{�b��1$��#�!��č!pQ�nP�'��<�"
�1<N��?�0�7�gyB-
�߲�X4�� �U�D蒉�y� �.@T�Teε
KR��D�շr
r���'08��7��*T �Q�-�:7���'��Xi�D0-$��T���<&�=��'Z8��VKZ�m4�`x�E�:�ʱA	�'�䁨�XS�L�b4O��C8j��'ؘ�$T_��{v.�Fp��@�';0,�d�93��Ӷسh^��A
�'FFD�ImeR�9���R\0�'4�̓���8&��̲$�U�`�h��'K�ʷ�V|~��Tj>�8���'���a��J;��� b4R4�	�'"�d��\&l��+��!`�Bq;�'�v�k&�[I�R=�m��`80�'�pb]����T�ڵ���s
�'0H�@ƎB�q� �	�
ޞY
�'bJ�j!�D%E�nY 3
1l��9�'�&]1��>3<EÒ�]#b��!
�'�f)xѤK3D� ����N#�4y��'[*���D �N�\t���A98g�`b�'�ر��N(ZH�1V��3�lt0	�'�,9�b�@��jr;(��'ɮ4C@*
�	�щ%���#�ea
�'=h h�M��T��#d�
�[l:��'��� e肪sJ���FH�jj�y�'O��(4+��v��8t�vX�
�'KJ��� c֬f�
}i��
�'Xu  ��WVx��D�n���
�'Gb�"��G6+Y��;D�H�7ǚA��'� :P��!U;�*�7!Xb�'ʬ�bq��&y�P�a��<"���'�r49�Hc���kA�?5OV�B�'�(�Cc�*ei��;!�Ŗ4p�	�'?��o��;�4s�e	0|��
�''^�! Z��� s�d��f�h�'��a�SGJ!0�i���>s �lp�'d��a���2�z����6Tm���
�'&捻K�,|؜��D��J̞�i
�'팄�B�;��,я5"���
�'�4 "c���d3�5�wK�*�R�a�'��Y#��;th�(�Y:l��� 
�'��a�� G{��遥Ǣxg�<J�'2��3E��F�>�A�K�Y�X9�'�)��k[�)b!	 �SD|0��'5�d��NZ�n���LG,F�=��'Ȃ��	�_�	s��ٸ&��)�'��9�eל{��Gi�gtD�
�'��C$%���up�P"
�'l��S��Ls&�:rDͧ$�����'�"�L�"� Q�kI�e�v���';Q	§@�sr�] !mH3QVd�'L�;E,^�
	t����_`�Α�	�'�t�Rc��cg�8��dW:�N���'����Z3L$�TH@)���
�'τ��!�*sܬq�BJ�+f�
��� 
�;򈋐MG@͋Ԏ\4���Y'"OҐ{6̏+������S/O����R"O̥ɤaD�N�,X�𮏑&�AX"O�Eöń2��e����6Ln9�"O2�覨�0���W#�"��(�"OF 3U�E����ŁM�:�LQ"O�	�����0$c��S�� $"Op=�禝bqP0+D
ѱO��S%"O��Y�%Y�d�pz�+Ձd�P�:�'BB�1��K�4�]0�Ƌ�H���S�'��)4dL�Qa0�x���{�*	�	�'�\���
�a=�X0�c�/	n����'u��Hǔ�8�"H��V&��m��'&4��&�ƢG4dI2�Ë<E��8	�'�ԳP�Ō����uB�-� �	�'<J�"��r�� E�#%re��'���@O��!�.e�&�1+L���'�n�;3�]�Q�B"B$�� �	�'ޠ��%<W���JI��s9�9j	�'麥A`+G�*~�p�'+h���	�'6��C�@4!�j���^��	�'���xEgǇK����^�\��'�DE��`�'�~݂�Dn��a�'NV��PG8�aS��]�vı�'�x� �!SJ2xJԪNP��0{	�'���iֻ9�ɸ�CC<N�f���'�H�ss
!V�Ev!�798�`�'2�Z2N��T�Z�镗��9��'�6E�4e�)q�8���f��8�'7�1�`f�8e���l\��f;
�'o���]X��W�L+CD�
�'������!X� ��N6���q
�'��iH�>M8�񃃊�.i45��'����ǔ�g�$���./�r�'t��%A#A��YBMI�S�І�xܒ@���]}��&�kr�ȓ.��#�,�7t8��bG��
5����:Rs��=p$ ��H�`t���j��!����}�@���l�'Zj���?86���'Z�X�ҥ�c�J�I�)��&34�ŠC*dKB�N0	���ȓ^Z T�#�Ճ7�`�As�،�J�b�=y!VF���m���L�'7vI@��G�����+!�,�X
�']��k��3D:�H�!�dª]�4P��}r�LρPI0��HP�K�:TF~�`P�w�>(3��_^P>I���۽�0=Aҫ?ߤla��ΉE�I���Fj-2FY��P��!!ʧT/Ρk��' ��	1/򔚶��j��h�<���� J>�ihJ� 9H��*G����TH�,��_�T{��;zLh�I�"O�qC"M?[�@C"F	%�~8P��X>w�����d�T�R��i�"|��T�l"p�.*��z��\8�1 ��.D�h"'-�h,Jy���<W���.w�$��U	O�����"H�!����F�ɻ~Pe���27�6�y��(.�N��D�]��=mA���,�b�T�T����7<�=��-�'_#&��E�@E؟�Z3M¹2�t
�`�&�6$k� (�6"96%i��uS$�)g�Q�@��i J|����65�p����!wP0��-!��>Pr"���l��)�0��K�|�!/ұ(H(!�r �2H������ӛ���
c�LY"#I+F�m*��ΰ�!�ֈ[�QA��ނppv�K��]>G��!5$��,
o��$Z��u��X�'[V {��j>`r�g� T�H�
ӓ _��ұK0j�P۶
�#VBH�RfJW�B�z��&�.F=��b!��%&a"��0:5�ɷh
2 ���vUҘ'�v�t]rr��W�κ<�!a/�	��g�B(��_Ѷ���
�g�!��
c'���
P'<�T��e�`�1t*I!:. bt��.ΝR��ә���Z�(�Ҵ;�뚠W��;�*���!�� <�S�-��M+D�HDO�_�4�[u��ذJԪt����DӠ0��F~��7��9�?[B�$z����0=�=�<�DM�]�٪��D�T	N���O$T��рB�J�LuI��'S^ݱt
�4@���s��F3횐�y��N��7��='�HPC����ඏDD����@�A�$ZTī"OL���hX4d��9zgfM#�1M�3vp0��.ޘ[׀
٦	9��	�d}2�&W�0`;��0��Лm��y©��]�D0�wCE8Lh�K�Gܿ�M3��&}n���-8�����[_�':�R2O��p���a��¹~J����g�f�bc�TeJ@a�e΀�5�����.�� dE�:u`Z�Cha�e��V4J!F@�7R�8�j��'T8�n�/���bdU�T��{�t��j�p�*&K;$r�����80�~B�I�6��Q�$� r� %S0!�)h>�TiQ�5�"3@"%S"7��N�O� �{�Hl�� 6D]H�s�%�Ne6�ȓV��]:C��f�6}�a�I�e)��mZ�k��H���Ɔo��8(�(M-��#?�
�5#ܬu��G��v����Pm�<���:B��R L�~l�4��!Eg�<�f�ܾR�N�{����@�:(�7A~�<�˒�B�@ȸ7DˬD�*�h�x�<��^�>dTa+�Q�J�ؓ�E��<�U��5m�D8r ǥ�$��D��{�<qB L����A�%u� [á�B�<��M����J;��P��Øi�<�/�3~�h���^8@�a�U.�\�<qK�4���V�Pp�+�Be�ȓ���[�х��H۳B�%.ˮ|�ȓ$���ˡ���e@҈(DU��5�ȓ|l6�	��8e�`y�֩�b�(���0���UAϚ��0�aF� l`Q�ȓ����Gٝ�P̉��G�&�Ȇ�P���0��D�����	�;��ȓY&n�@v&B:�������6}$���ȓ3���'��U��D�ƉW1x82	�ȓ\@��)VKֿ �^!�pG�4�f�ȓy�r�gN5�2P�vD�	+����ȓfo�(A�r��0��nI�}����v��*���2UrP0`�I��-�41��4w���.TȽ1����t�fX��gR=��(^���c3��}ºL��.��}�C��	B;\foS	P̬%��
��RWN@�ej�����R�i��H?��яL$>�4���K�y��H�ȓIB6�Q/��9���B��ݝFJ|��9P��s�ĳ}����G�	\U�ȓ���"�"���B�P��^�M�.I�ȓ_E8�� �T��ۓ)�m@݇���[���:JL�se,�.#����c&��:��)G*d���*UD��ȓF��}��I��[�xeS�f*L�z؆ȓdu�}9ᢗz�L�z%
��I�����3�&�Q���v�壶邠z����ȓ3\�9ɁH��^�FԼ6� a�ȓ]���
��ԀiF�l"��U"c�)�ȓjaਡt�L6$�ȁ'k
*V>��Bd�Ġs�Lu�iq�*Y�`���ջ��Q�@�!���$KF�ȓc𡹔FM�>�8�Z��h}�A�ȓ	2�2�k
e�
�"�NK=H��ȓ-�&IP,@�Z�b,� ���p���Io�q��ԔHE@���l�&ȓ��B��L��pe qE�^��T�=���^?_"*e���*'��Q�/X�� Q����#̕/x�V�Ap�#5H@B䉓>>Q��b�_�8E:�"�%QB�	�&W��BWc�;	�QG圅:�$B�)� ���̄�k��Ņ�99���"OD�Q�� P
�1$���
jP�"O
x��E�rX��q�,_����"O(,I�5n����F��<-��c�"O69�POG�^t������L�QR#"Oȋ+ڭ���1	ңV�8�p�"O\yA�d���4��Λ+z��"O(�Yg��y]&�1!��k�`�U"O4��@� =Ir�gF[#c�D��"O,��p�S8@7��H�O!�m�b"Od\�+]�RIҐ�I�C���+B"O,���l�>hy�u	��YUZ�(�6"O��(���	�UԏyK�ڲ"O U���6bbzm�����/B�Y��"O�<�����?�$���bY�1RDm��"O�Mb�ʟ4
�`�i�Ⱦ(�@١"OJ}�I�ZA �0�չ�"O�Pb �"� \��`ϵb��)e"O���"b׉ZBh����0j<`KA"O@��b@����ũ7��?s�d��&"O 8� L�+F�P��'�>(�zt*""O4]�K=�Zʅ&\1�p;v"OҔ��D rB�k�k
��A�"O�|�!�r H��a���&��T"O��c�_t벍h�i�+iuV�(B"O�=ap�S�F� ��탬:vD=s�"O�5�®9s
0
!*��?��Z�"O���&�O9���@H�,{ �G"OrA  )џg�X�F��I�,p��"O�l �o�.g�("��6]����S"O��Z�Ɂ s��yF��6��f"OP�p��H,�(#��Nf��e��"OX��Wϊ=�҉)�d�9�$��"O\鑂�5Ǹx�b�	�D֚hQ�"O~��E�4�8��g�P���R"O����%�G���W�òV��""O�u�q	#1�V���/%&9��"O�p�T̘%��7���J��I��"O��+���U�"bu �)�$y�"Ox�CmS�~>jU�UiյF�����"Of�� �X�"��P!�gς.�z�j"OR�ɳ�W8\�0GG��v�ը�"O�L3#��K��rk��Wx��u"O��`��L#�q�$+ʔlA"O��d
�� f�i5L�h�$�2"O�("����h�>�V*��b����"O�M+ぎ�A����ݨ<LDlS�"OrDI0��\cʹh�C�;�B���"Oh�8�ׁ�t]�`�E�Jͮ�0'"O|��bA�qԀ�v��8�c7"OL�0�ا�P� U�1��T�"OF��g�S.w*XuSw���q���"OLu�5�E�0nrx�ړBhj���"O���0���Ed<5�ץ��Z��s�"O���@�@q�}Ҫ�"yr�Ip"O�(��e�d~���Ơ�D��|@�"OZA��)}a�f��=��P˦k��!���X(A҃L>*�80���)_!�����D���K�μ�σ >^!������Є'r�A�o+Pl!�$�YC�1se�u^|�B䣜�1�!򤟻:�4L�Z3^R>�H7�Y�8�!�DJ�gB��VA'P�8ʅgJ/�!�dÙx�0��ˉ<v9���f�>I}!�� �u�Y�U�X8�6Y��Q�g"O��I��g��a��5^nTIp"O�ٓ��k��@���1�p� "OPK�ܹwT����K#N��2"O��@H�aGD�@�{J>���"O�`\�L�M���+,�5˱"OU��/�B�Z iHn(,�*�"OP����P�p`\l(��=��`"O^<�Q�f�H���S�G�"Ԩb"O&��ч�a3��;ԎL7��q��"O�����2)��4�oФ��@�"O�DTm�(~pO]8�X�"O��[C 
��f]3 Hĝ��;S"O���@�cr����x�|-��"O�(pO�H��(�!Ŝ�S"O�)�r#�6��(1� #D[h̚"O`8* �r�3��ӽ'n ʦ"O1�����$�����ΐ���+B"O��K�LD./sP��6�ǎ:�)�"O�XЀ�P��5�2Mš$. ��d"O�0i�J�6�v9D��(D�p��"O4-�
�QB��P���_�q�u"O��{�*�20h�F�Z3���J$"Oh����
첔��f�>45�R&"O�l�v��=
���%eGV
X�8�"O �CUG'���f�E�d�	�"OJ���n��1,��S�A�Q�KU"O�E�*�#KQ�i��n�1� �(F"O���bܶd�$��ϐ�o���"O����$@��L T�G�UF���"O衉͂n���H�f=���"O��`a�r�Ԋ%��N9ZqJ%"O$Yb'O�
0��a�FJJ�&6�8�"O������4T|.��E��!I��%��"OLT����`��#�Z���"O�5Z�Q�p���(�g� �(d"O�lô-ހ=:�n�)�ؤ2�"O�}rF�Ӫl��a�m�e��u�`"O.)��
[Z�(F
Z�m�r�c"O���3���Y��Q���8�b�"O�d�5�!?6���F~ ���"O�i���"(R��&`�;IfM��"O���A�ЍR��y�cL�7Zs��v"O0�:3��H���6��
s��t�"O�����Z�(V4�Y�e�	��@:�"O��@͌\�Ф��dM g�s��|��)�Shf�Yi恙�;f�(�T�� Sv*B�	�R
t��D��) XT��!;/CB�I����5l�G��<s�%
�yF@B��8k�qpp �<.ܸb�M�3��C�:5~L��"Ѣe�Ɣs�
�\P�C䉩x���p�K��~���L�'��C�	:%�F䣧BQbo$��#�M2[�C�	�r�r�c�%Ӏn"!���J���C�I# ��X�+Ё[QZ�H!��6C�	A�иh��F,,�N�B`��*y�C��=z�������,!�l:o�C�7y�,���D%D�lEB�� M�NC���(�7��&�D�`b�C���He@���$g�|5�֦�bݠB�	%\b�8 �Z�(fp�ʴ"@8zBC�ɋG�eh��8B� ��E�J<C�IM1
�d�M�,��K��G�B�	�rw&�����{h�S�8��B�)� �2��A@���,݉<��@��"O�Us$�S�&P��b5,�{��YE"O�Y�P%ȯx��x���-"\��1"ON$�Ս�5Gi!�j�l'$�#"Ob��I��"W���]�p��"O(�6΃:ɠ�[Qˈ�uY��"O4��� l DPz%ۗ>FI�"O���-K��董�e��;@"O�\B���	_���8��֓P����"ON�{� Y�R��eɲk&.?�@ʗ"OR�
S.9/h,�%�uͲ9��"O���C,F���y�H���j�CV"O6��$"\�|8zg�K�r��c"O2��F��2Y"4P��:jr��"O�طC�j�X�a���$m~�hg"O8MC��V]�k'o�|a��"O��X���I
t@��Y#'�q��"OV�"n��t"X�{�� >Ґg"O�\�憈1q���!C�,:NM�"O� �'�<�������F�r�X�"O�|�L�b��Y��� Q���"O�Xb#	�7G�
����)�=��"O`�`��N٘��B�/3e��0%"O\��g�Z�H��y�Ĳ@"O���BF��3�6��Z�"O°�`m��I��T���N�̚�P�"O0����+��=��_'.V���"O�:��ч-��e��:;&(��"O�(���OxS�Z�g�0Ӷ"O�̀n�+fB͘��3S�&�2"On�Ba	ح���Ps�s����Q"O�xq�	"Nu��t� ���c�"O��D�
0z�5����}HX�"OP�� �%+$��5I}:�ڵ"Od,�V!�\�:�I�"��g�X�H�"OT���T� ��!�ҧ4F��@"O�p��.eX��'��#o��t"O��ې�3�-��z2yZ "Oƀ�R*G0Ӫ1
��۳!kԈR"OH ���6�������:2"O�i��bݿ/�84�PIV�|��Z�"Ot�(�^Z����g�ޠM,T�"O�HB�yh�HBP�@��Ś"OFiq��h'l�`D��&��}��"OpUR��q��]!�˩L�x��G"O�1��@3uϰ��
��kB�i��"OfI�ӇN�)�D���/Zz5A�"O�ő�i�Ch�``fDۄ{��	2"O~��a�Dy8��L��`��w"O����7�qyG�O
z��ua�"O������W$�H�b
m�TUk�"O�8HGV5P��1�C��lH�c"Or-�C)Q�]:��+H	�R"O��0
s0�0�h��d��ٻ�"O �PbI>ڂ����ï5��=�a"O���	f�r���f�6_��h+�"O�i��K�(����D��qʱ�"OTPQ���/hh��U�d�"�v"O� �Ǚ���*��],t��0��"O�{օq����Ǟ'YJt�E"O2�A�� z��t��+71�P"O�y��#]�U�lQ9EN�#0�4d"Oh$�FƄ/M�DY(���]�K�"O���c�:Q���;�l>c�4 �"O� P��%D=n�!@U��.�H�C"O��1���[@��rSI�7QrnU0�*Oj�s4�L�,N&Aң�˘57na�
�'��|��≼D�ؑ�u��/><���'�~XH/��x2R����&6�zի�'G��X�hT�6�a��K�&�@4��'�Н�nJ�',L��+w�p�A0"O���'+Җ&�:m����63Ƅ�"O8�ح}�LD�
�qQJ��R"OV��G�:���qh�4,*@d"O��BѤ,�"��Ȕх�u!��9��  �)�m�I��D�1�!�$ؕ�DZ��\+Q\mx��yq�
�'��}"g�
�M6̅��Z)��a�
�'ӌ�J3kËV
!�%e�дj
�'Φ���:oP���tF�m�Q3
�'k���Oˎ^�Z�a���]#(t��'v�Ep���dh �%��Zp��'�ΜQ��K�J�t��L� �'(@9S��!XS�L@�bK�X�2-�'�>�PU��-Ði�sb�g9P���'T�([��ςTQX �J�9X!PH�'�J�2�5 l�{$�* �N�s�'�@�����,� �JH*	���b�'��uK!��!B��չ|0h��
�'!���3"!t�4Q�W+Ky�� �	�'ی� ���C< �J��	&�
�'��t�2�4����c�y[ؘ�
�'H<���G�
8��#C�b7�ə	�'�E��+����hz���0�*9�'�v�X��qx�Iր$���P�'v*��B�5T~����%Y�A��'���Q���~E,���	K��0�b�'����cEox�K�n����H��'�P�����p�!!��E�4��'��|��#ߐ~j�y��J�5�����'~�%�C����˅�(.���'�p�Y�]e��*�L�r����'+�+B^�&@hБ���e��
�'`�����+D�$�s�G&.;$�2	�'=��gj]�[���8�(�,�*��	�'fr0��/��7��-�+#@�m�	�'�\q:f�\N�XXp�J�.�{	�'&��p�\�&ٛ���GB����'�* ���܀]�Q������I�'�p��4Kl����N]�Y|h	�'	�t3�!L�FmX�b��T� X		�'�ZekR�߼J���#�Y�J`�y�'k�D� ���S̀�>i��b�'�P1�塀4ږ�(C�Q/�Zm��'���R���7])H(y�B��
�'ڀ��f���ABB�n�ج��'peb!�A�+�t\��kժj]��'K��Kï�=Y7䭰 A�6���'x����"����h�I��`u��'8u��ᇔ9 �}؇��R��!Y�'o\�+p�D
W
]�G���I��ձ�'|�q7̕rs`*��]�M28�2�'�jx8T�V�<���U�[�=r���'��Ր��H���1����BC�0�
�'�B;0.M�,wN<K�K�+��B	�'�.Qy`$M	t8�|8Wk�./-Fu�'��q��L�k��䨕��*A�:�'�B����)�č����1(p��+
��� ʉ8� � �䙢I�8FJ [�"O�4�dA��D�q*\=�Ւ@"O�9�U�"��h���2�-@�"O���mX�i���i&�T	aP�q��"O<4ГC����P ��}(�Q"Ojz��?C��t�A$Z��$"O��� �N�Hh�`YB��"O�麴�ӵ�F�!�7E�&,�"OBd
�J>q���GbU�vm*�"O^��6�f�L�c�N��`�iw"Oj1 ���i�� �Q�p��T"O��fAG�ZL��m�i��i��"O8!X�n Op@�Ѭ����,��"Oά�쌼g�
�Ic"Nn�V�{�"OdI��F�|L�\���� ykj�g"O�H��O"�248r��<e��d"OT���ʓ"f�Rf�˽ s
9�C"O�c�_��8qzb��;+�4<��"O<��r���%���y��"OfHB�d����Y���Z�:ӗ"O�IԠ>m V�9!H[�7����B"ORS�l����g�^���V"O. #��Y#.��00��,U�d�7"O�u�r  �ͫ���0lE��"OJ�"�!՞(��Q��.·y�>��$"O�<��!�b�h��E΍&���@�"O��"ˆ 3�� GL���0��D"O��h�	�&�m�U�X^ߴ��v"O$�b��{`��.J8�D���"O9S� "�q���$^���b"O�bq�Ӏ\��U��
ˠ?�4�c"O�A�%�.e\�Q�a@�>+�q"t"O�@Z`�� Dfz� ��C����"O�}�7�Ռw`�`��@�~Y��"O�!pF_!	P����,�9�!	�!�Dȹq��9��_W� ��q O�6�!�2Ud��Qb^� �Z6`��P�!�D�z&$��P�Kpn��@��!�D\Z���#����5[��b"N6m!�$�O�t�T�xQh�7/��lo!�䂛@0��)8�S�mM�Vc!�,��Y@�Ƞ.*@��w�H]6!�DǙil����;VŒL;!�d�(�L��qk�>8ֱ��ۜX�!�DI�`��h�2씢W�VIp�G�/*�!��2Yg�)�a�>�� ̄<'�!��7�����)��E�s�B�7z!�[�K޼���ɕiҠ�GT�y!��ϿB�8w���o� ��aEÇIp!��)#�d�p�Ǧ8e�*����f:!��Ϸ+�*e�N�z-�Y)Q'\&6!�$	uͲ���nB�I��LP2@�77!�ԍ���3 ��P(�Xe/D�+!��K�_J(p	c,�S�ؑSD�L�!��7Tyk��h��b�Y��!�DH�j<�'�ىEq�#k�!�XO���IO���D5Z�S�*!�ص7�����1�P�Qw�r!!��S�@|�����mA-�1!�D�u��Η5U� Z��́N!�Ď�Um�$��"5.;�D��2]!�dȱA�R�rT�P162�[��"B!��X�uvQ;�j�b�RȲ7�	]=!�dY/7ٻ���4�R	#�C�=I!�� �4:��� JQ�A8Z���"O�QY0�N6=E�n�垼�0"O�����(�
w
͸�< "ON�
!CV(�֬çH��x�`��"O�9��Ȑ�MeƩ�-�Ȝc�"OH�Nɬ{$��LI�1�-2�"O��#��1�$��`̒;�h�%"O$��Å�b��vJ�5ͼ�(�"O�!�2G����Q*v��	N� "O�-�������I�ǔ��Y7"O~�aI�%C�Y�%T0+�DU��"O�dzBh�)|&��fO@&�8�T"Ox8��!��@�]����;~�|�B�"O���Ԉ�i�8|Ar'O�C�(��"O�1b�Ėuyڡ����0n��"O�Dr%)X�L	2��
��JTcQ"O�BrW�1re��ֵp�8���"Ob�x��SS�pD �ǲF���K�"O�A��$���z�gŠ�T-"q"ON!�p�^+Z��� >�k "OZ�B���6� $��/��ބ`�'���B���)ָ�� ǽ 8xs�'d"�pRX�c2�����f�Mr�'"J`�&+Nn�����,��	s�'i���;D5��QǦ�!�R$[�'�Yb�)
�Xr�y���;9�iA�'+�e!0d̡_�:es��* ���z�')�ua嬑  Y��`�+�q,\l��'�>���lp��mS��E0}��A�'s�5�>R%���U(ִyC�i��'�yj!�q��q���}�8���'�����.Q48ƪU�&x�'��0��+��j��E �9z�&!r�'��e(I��d��ё�طlϴ!y�'f ś�J�E?:5i��1O!q�'�Dljf��� �dز)z�Q@�'~���B��\#��Ӭ!]t|��'��X+!��Yf$��/�V�|	�'�8�yV��R����8m� ��'��Lh4���p)��PƓ b���'��h����(���#a�E*eФ8�
�'��͐%d�=Y��-�f, 
�'g�uqA��Ei�H���XXϖ��'���0�v�eP��5V�HQ#	�'�.0�2k͸MeH�kc�ՓP��̸�'Md!��4,�p���5r���'c�yH�C_�@҃3m<%��'����BߤO��	�«�';Wtq�'Q�Z�ȑ�%�2���D/1d��'C��JQh׳H%�R�@J����q�'�&�s� q��Ta�,(���'*
q��-\�sq�DcݜJ�a3�'�Xp��0_s�-� S�Bv�(��'�Z��ʐ�`���ƕ�8�`���''�qï�u��x%�W�,t�(�'���φ��J��@��p�8�'K"���(M��l�1�_�v��L��'Z�d�&�{�>�yD� o�>��	�'1P�j�.̽hh1��,W4z\�m��'h�h�a�6�`X�1�o�����'}�h�R�S'��h����~YDI�'�*�Ȅ]�$�����:{PHP�'"�H��f��0u����㑣 `�1��'�.� F�+9�#�"�f7������ �D���5T���z�&�"O���Ta�r�0كA�Q^��uS�"O�л7L�h���I�X�\p�G"O����N��iS޴�vm��>o���"O6 h振{��`qA-�v�U�����L '艚\����'��tW?ib2d	u���:��\�9�>y�g �&\^h}����?��tJ>��淀i�N<)����*@i<�;��a#��� B�Ҽ�D�]�V�j"=�%�l���e�M�G^�k!�A�w[�	��+���B1�P�0h���8"L-Gx�c���?���I���'���<L*�����75#0��B�.@dt���������A��b%yņ�� �x�Õ�Dx�=������i@ݴ�M���̇F�(����!wB�w@X]?)�#[�)������?�+�P�{���O6��a��x�2G��:���@uY?K���Ȳ΃^�@�gG a����k���џbʧ�rXc�6<�0�Ƽ0�����P����4coa��^W,rҌ�(k`�7g��X���|��n�^�B��So�"$�)��(�Ŧ�Ѕ(�O�@l�/�M���눟���U�W�&Q9���-Tl�ad���~2�'���UX��"�"w��A�oÌ=��t�`2��McѲi�'��&bK��@��@0yqEH�l�<`2��?��ꍀiBz�A��?A���?9�U?�n�4�8e�$�C7|�J��K�n��8@�S+xNj���%
0f�t��u�Ǘ��b+%�B]3���
���er��sqK�/��`�L\�P�'Te��&�<�<��ꈨ���
>�I��A>ZF�����gy�n��A��ß���4J���gy�!f�`�JcP�ʰAU/'�N��1�׈!P�ȓA�.�1�M"^>x��G�Ħ8��e�>�mZO�Il��T�x��˕�G~eKV�ѕr=e��YI ȫ���$�	�$��/.~}�IƟ�	mq��mڧX�J�B��=_�f��b.��c"A��VJf}���OF���OaBFN�|l��ī�ǡ�vsΑ�%*��G���Bb,Iߦ��3��9"������߳�U�4�M�fP>x���1����(I�O`���O����Ӧ�yDi�>NA�hZï�|s��g1D�����	0����!%�5.���n��ߴDV��V�hBg�%�Mk���?��Č{Ra]�Q�`k�%$��VN�2z¡�	��	�D��	�!��gxV �MS��Hp��8���+���Tkp�=1⾰k�鉋Z�L��gFl$r�9r�P�E3 ��Տ�j��
W��	r_FHR�J?�VႦG1\��0�I͟ �ܴ�?i��T�	�-L:]��r�Ŗ}���5IUݟ��?�O��O@ٳ�_2W�P)�g�
l����'՞7�����o��Ep�2���/N)�e�^"*����
ٴ�?����I��0ud�D�O�7�E�F��%�X��JDτ�#^@(v��e�w��h�0=)�i�<���Sg���OkL]/A�!Ǩ�;��#�.5�f��	���d
,b����4Ob�`��ԸX�1�kL"ZT�rт'#(��]Vn���>�?��E��#|n�V�����ʙ0>.���.S�Lߞ�	ڟ�E{��d�>mۚ Z�"O��8�Aǉ��FQ�T �4yݛ6�|2_?�� ��!I�2-Kqh-@��sɅ����Od���1 8  �   c   Ĵ���	��Z��w�D�8,��(3��H��R�
O�ظ2a$?����`��4h�vGޒ?M���Am�`�8���7>�-��lӦ�lZ%�?��'�V˧��mZj~�ڹ���G��B:���F)^fPV��N<!��=ζP�H>����a��d@8Z�0tRb�;����eh�	:*�F���
D;t]���x׌�F���/O����*YN�N�@�/�����&0�r$),O���>
!f,ʥ���W��ɕs`�\a$��QMؐ���T�q`�ͻ:��}�UU�\�*�4����A�<1���LS�o�5
�|�Zс�9�@�S� ̋N��M�_�0���{�Q�L��|�F,^�����k!�5d �y2��S�'s�AExrlNqR�SҠɂJ�DP��яEo�"<�28���lS������|w�B'/gA�O���� "ϸ'��ab"H\%\��`5oʹON]ڴ3L�"<ipf6�!0͒���Jv�����'"y�%,�S�Ǿ"<1�'?a2�Y�#��(@̑�_��0��Qy���N�'���?	����V�^Y�B�·cb"���_��#<��,,Ђ��G+*�	��c��Bl���P�\9K1O���d��A�I�_�L��)��hZ�!�����'��"<��$ �e�}BCJQ�h$�A��+��*~��矬�]�$�k�a̧#t��shk�A@s`� �԰���]R�	��M�<�OՂD����<Q���G�Oȑx"�2F�bբ&�<�viy��'2C>-�6�)�ԟj�Ey\0J���x�!�`�|����y���h d  �^k���@�:��D��d����ݾ<��(Z�-�n�YF��*����C��4�џ�: $2,<P�S�O�0�&�1�۹���D;0���F~"��k�Ľ`�O \�e e���c3�\�p{`{���3���3o�w����O��qР�J�@��`Cʑ�3
|�1�b/0�9G���ŒWĵiu P.�P�Jd/��䕀C[�X"��?om���0�Y*��̆B H�A`_��!��G"�HJ�G9�`�һ=n$��A�"�򤂸I���1�/��$��A)Č�FDF�p�ƭ8o]CB�2dܧB.(yʒE�3�8!zt�W�z�q��mR&/^HL �'�*��� �5ɈE�L�yu\l	Ó���`���:b��'˜ii�͖E�JP�թ�0@��T��'�$TtK��gi5P   �
  �  o  �   �)  E3  �9  �?  iF  �L  pT  �[  �a  6h  yn  �t  �z  C�  7�   `� u�	����Zv)C�'ll\�0BFz+��D:}"a��6��ԫ�7O~�#�<O��S�eŲg�ء�e��b@��ۗ���ǧ�ũM�3v�9;�i\`\z�Hdݙ�R���?�W���?��B$B�6���C��_�`��P>J��V�5�\d1���6�Z�����u��?<���m�V��"�|bQ�pˀ�F�����X�x~�梁�����$
Ops ��M+�I��?����?i��?�Le�Nh�5,Y���x��-y?ʭS� [	Q;lX����?Q�'�1L��<���?�T$��k��IZBI[�e�Q
��?���?�����OH�e��e���?���^O�č��u���`E�	�HO�0ړ�M[��P�J̓���(Y���𧊎'����<���$�,��8�O Ġr#
��X����s$<�V�'8B�'���'��I��p�O��A�k>�m�'�"W�~t���՟s�oy��l��M�$�ijOxӂAnڶ�M�`�iN<���1�dQ�U#�/�<���gk 7��O�2��;i���DG�!b�I���OvD��3W�ͺӃ9p���2�ѳ0�F9CAK̬x7��3���/ ۪8o��M��i���ޟY��-�$Q�%� ���h$@ǀN��Ғ�id�S 	W�ElP�߻_Ұ�mڌ> @�Q����u��4ڛ����W-�31Ɓ�F����B46 (U' ��cyӆ-o���M���\����D�Mʖy0�`B�r�fr&lQ0i�p�����J`{��� K����A����v�n4n��a���T�ڰF�h乕�5FPk-SS�e�pf�r� 0�!ɏTWB7m<�M����9�~ A2��a����6�ɻ���s�@n�j����%k����I^��?��U,88r�iiR��p�'N>��CԳ{���*�� !F�p��S�'B(A���'�i���M�t"R��Y)�O`}�2j�)guP�����FX�U�'Ȏ�nZ�m�"!���m}b@O�qlF���Ox
�˧��1�0<A�ٟD��}~,�?5
��5�<:�NJG�-�?q+O�=�}��钘!5�L��kF���DnJ��\s�	Zh�7�M�0�^Y	&�E�v��z�}��IG�T0��[�(��]�
�#��"�]�^!��"zN�{��B�A�>��R��\c& ��T�d Q��Z6\0�-�,',���$���Ahh�;��i��U��7W��Ht@O��TQ�OɅȓH\�8�[X}sa+������M��?���?���?����?����{�f�L�-�^����pQ&��n<Ui�雨W���"��$E�!�/����F7�ēN������խ[�|03� <0dK��Y�Q��CŚ#��$Xq�W�N�&uZ-�h(�q�j��?M����a�;5�\q ����6-�]y��?	�'���|�)�
�&����6�:���%�j	�'�b�'�I���i��J+�Iٶ%V�,���F'6�`e��m�R"�'U����d�|�����i�m<J���A����
K�#h��y6�����r��!�B&�`P��h$<f!�D�S���Y�.
�L�\��!G�Ec!�$��hY��S�`'��Ũ?P���9:�*�9$&�7�L�����yB!�4��!��B���a�! ��<����?1���?iC�J|�h��*T5ؔm�b��&�?A��gڍ0��?	��|N��� ��ȡ�R��y'E�fD����I�C,H����K��0<!�,��S"D�-}���C��`�h%(�Nؘ&���1�^!.>�8���T;a��l��Ml�˟4P�g�3z�P����Ժy�)j��͟��	ϟ��	�P$?��<����0mbL��C���Q�5*A��<��	��M���֖4~8
�R�88�Ԧ	Q�r7-?�	Ӧ]0���Z��Z�ŶS�42�!܎��b#I(�y��S Q-��!�.�"(�m�
�y���%Ԇ�;���N>�`0�y����P��2w�J�șr'�=�y£܆"\|i����ؒ$�@D�*�y��ѿ;B���G�N�&��hv-�>3˛�'�r�'s��J�~z�'-2�'$g�\��B�JB��8<(�ð�a%{�H6{t6��Dw�T����|����7o��I`��J(^�q�䈲;�x0 �5��M�`.X�����)1<�C���e�"��/|��<�t�şP�Ƒ����?������p�d!\�z���_~0�c�'l$�P�i�)�L�;�DQM 	�,OX)nڵ�MM>�'��,O���Ŏ"�:!a	��!
μi�cV-N �BӉ�O��$�OF���⺻���?I�O��1� ˙����Ћȏb|:��f���xR/�� ת(�pϞ�٬�:�오K(ͣ�'Т(��� �>O�) ��W�V�`@�X��?���'a'Վ��s2�Ey��P�'^֡�@�@�XS���U�؆/j�L>��i^�'�-[#l�~��� �X��2��p�ι<Tް����?�#	��?I����B�<^N ��+5�p�i�� 褹�8m��Y�16V��("�\�\�ÄG��d�H�pGm�8�M�K�nPp�S��ʠ��AべC���F�\��OFT1��':r��h�'��A�>���ޮ�x�Q�/��>�O�Hf��
���KQ��J�f��f�'����Ųba԰q���A��m#�n�/_��W�t��"���L��˟�O�A�5�'q�pj���9zjA��M���pu�'k�g�����J�	t�>�kd��Jz���'��)7���8C�^b
�{Ɬ_q�ɹ��S��Y$K�ԁ�@ߏ"`3Yw���`��,��"��2gǕ��͘ _ ��$Nk?)��h��o;>}����r;"������C�Ɉ\��z�ɏ\b.(�4�_,{��?٤��*|�cM�o���Z#ۨm�z���Ov���O��3��^���O�d�Ov�3�es��j�|�S�++��0,_-q*E�E��%���Q�#�Ӫ��f�F�C�`H�Xu�W��$J|��Q5�\$"a��(¯Y�e$���$��'RJ���i���$�x`�cb�X�x1Ȕ�؉6�2���z�'"�I�i�1�I�k٢�Bw��:���Eh��p^��H��"ߺ
�@��'ӆ"=ͧ�?�/O��p��8SN �"b��7,e���Eʝ_l�!KF�O0���O��D���O�瓀h�����8.�]�5��U���eE��,���F׮lS��+��3��O���3�B�]�.!*�d�T<xu�j�8���?n�@�ۼ�XlZަq���p�. 
���R�^`)��	7#��D���'�B��D�'?�H���֒Qw��R��D!=HФc�'��QĥEXc8]�d�
�1[�hL>��ib2Y� 8%����i�O.ah6��dqeY��/1UH�s��O���B%����O�S"tPW �6!�LBX�Q���y ��)�$a6&NR���C����O(�b���!��V#�:��<���00f����f�I���?�>�n妙�2	��H�In~���!��R�&U�&��<Ӑ�����0>Q�8
��`��fNT8pk�H��p��:�`�g��(u:�Qh 7,9��Ay���I��'V�[>�+R��ǟ P1�Y4o�)f��p�T1
�����ɝJ�P5s�,Ŏ"���1��_w �Q�۟��-kp��	\�#B�����w���D,?���A�n�:�R5G��00� /P=,��z���-�n0��-�G��y��N��tҚ,rҔ����'D���<�F�[�,R�U�cm��c880c��UL�<��:�P={��z��1��N�'��}�Tg^0W�H%�b�
Ɣy!w(�M��?��*�t��!�C>�?9��?!��ygi^�x�ݢR�Ԁ�a
K�3�m#4��%�ҡ�B�-�lTB��D� �D�:ٺ�$$0*��R`������*B'�� x�c0�+?ƴIp�	�r�=8��� L2l.���2B���#?�#ǟ��Ib�'����`
Ə2�~�AU����b�"O���2hđ��h2�N�7�B�Z�\y��4���d3?�Q"C���@rr�;Laz4�Q�jy�&.�p>�A�`�r�����3L��ʦ�A�<A��/rp�����˭�M��G�a�<9G��p`jʣΦ���Jw�<a7�ϴ0]BQ+��U�bL�6�o�<!�G�m��5�b�n�(��B@x��P$�����͔:�T����,���*��<D��quo�g������G��5�¦%D�qL��t���+Ţy��mXV�"D���EK�,d��K�5"���F�.D��x����k�<���-�jA|�r��,D�<�`
	+F�H�+L�
o���R�%�i�|�G�ĈO�f��:1L��5�f�P�y�nXi�KD9Q�7.�</!�d4��5�d/{�Ճ� H!��3f':8`1��]����Kl!�^;?���O�w�lw�YK�<��HM�a���+Tg�b�����ğh�n2�S�O%`�ĕ�v��3A�]C��
0"O8� �KU3I- ��p�\G(R�ؔ"O�p��'�O3*��7cگ
|�2"O������NT��Ќ�"#n���"OP�ҋ�}]ȸ��K_���t"O�ذPGZf��]�A 1���S�^�P၊7�OH��T(�����'�l0�9�"O� *1�VjO\#�m���C7���c"O����b�T��gL��;V� ��"O���$���D�y��,^�u�"O���gA�s8�x�J_"��S��'�!��'D@ 
�)��K�=!�c�j��<��'v�܃�oô>�&����f<��3�'�|�tf�%^�z�{ 
� V,�3�'`	c1JI�bv��*���SL\i��'�
y+`h�0aQ A	��:#�5�
�'����"y�4,��M�����dؕ\Q?�I&�"D8��R\�(F|�'8D�(HT&Z�c^�0bXT�N�˄B3D�|�@A��#�4be`J�F�l4�K#D���bҋgj�|�ь"iR��� D����Nz�H�h3鋔?RڀrTN>D�l�JD�h;�ɽ�-�G�O�MZ��)�'3n(�`�02�z�ڦ�B�7Ff	��'���Q�,I�Di���-Zd��'��� �h҉$:�a`�#q���'g�i�G%ۜ#��DwG�� �C�'΢mA"�o�T�v��B46Y�'��I���	r�2� !��;�n�.O61��'���[�ߦ3��bE���8ƌ��'6x僐�)����7a)��
�'I�<) �Q�V)"$��a�(��	�'7L��ԏB5y��(�-]"!�	�'�F��,۱. x�4k�4O>(3�0�����?��" ��G3�C�NԠqⰇȓ��Y0+N�L�d��K�x��Y��(���*�J�O�
W"������J?6a1'��o��	2�
��3�@|��mĭ�F`B�j�����;X��4�ȓi�HU�V��!0 ���<��G{�������u�ԇp\>	���ԃ0��q"O&��C��� �8" �?�:�'"O�� ��Ւ�Œ�Oڣ�|Q��"O�U��[�3<T ���Q����"OFYb''�v�h*3�]�?���q"O��"�&u�\2�Ĉ1P�0-�'�'�̐y���������*Y'Z5`a�E#i$�݇�v�3u�C�6��� ŘN�$�ȓ�-�0�F'qJ��c�iU����ȓ� )x��2+��#�!�n-��D���gZ�V�nXD��ՅȓM�����$8��XRÙ�kG2��'o!��a�6y�,;���hQ�5����o���yBN5"Z21@t�|���ȓV1z��@�ړx8�+��;z����ȓR`���W����L�ʴ��)��d;A�@*Qn�Ł� `@��ɻ��ɔ ���x&jK14=�Xqת��w~C�	?Cn0E9��8P���)f�߹ �B䉎�pI��K��P��BrΗ���C��(f_�y33@��I�g)B,[8�B�)i/ �!` 1�А*�Δ��B䉲K�<�#A�i9r乑BR�n=d�=iVL�O�4�� lޡZ9�qa���H�H}��'u��R���m~����42#4*�'+�� g5Y�900h؀'U��	�'U�����?^q�瀕 st R
�'j ��"gA� �����7CI��@�'Y���N�V: *w�K�o�n����!cIFx���W�@t�"c)\�KS���� M�tB�ɴ0}���V��5B�0�0��:�TB�)� ��&oJ0д��e��@�j�i�"O�����'c]bX7��]���"O^�B��	2�^�������1�e"O4pqDO��8�t� �)�B�gY�D(�G<�O���uI� 
�6D�o*5�U�"O�#O�~CF̡ Α{b% �"O1ZѩSe��<��,޺F)�"OB����&"��颦��s䒌hC"O�uK�A��o ��Ӧ�Z���'>:���'�0�O��*�����	�NT�h��'��h[V�ƐgI(9څbԄF?��'ಽ��3I�\h&��'@B��
�'V���w
(�*�2")"B@��'B���a��>}�6�(�-ߦu�<r�'�81`$�ߠ+�Uac�X�HI2��$�1�Q?�a�!�b�N����Ź�J� B"<D�4ʴJL	�ŅM�e�u�5D��;b-�0_�D�'�lH�BI)D� � �W�Ĩ�K�E��H� �u�,D�TJ���v˓�

H��`�&�,D�\��fN?@����኉C��8Q�#�O	�C�)�9mX�b*)\5B��Z�&�Q��'��xv��5VW2Uɠ�׵y����'�~�Aψ*���3%䘳!��\��'0~P� a^�< �������'5��is��;E��z͂6Z�j�K
�'�&���E�sN
� �]-<��u�.O0��W�'����(Gx�L�z��S.���q�'H�8�2Ə�NXX����4}��' �咐.ϕ.��9��3^l�e��'rp�i%�P�.𪴠�'�@�{�'V�Z��Nꄭ���U -��Q�_�fq�^S��b�5[$P��E��Dx��|�$�J�4���8��տ!�����3<I��aT�p_P��u�`k�4���m��HB&�-���ĨJ�D��ȓ�t�ǭN-D��I��O����M�ȓ:�:=s����"Z�Ϯ=@jF{�G���ȰI�b[Wr��@�U���lk�"OB��Ў�f�t�h*�x�9p"OdzBE\)_�i1��)<@�zG"O8�h��
D5�H#��,E:���F"O 0z5m73l^kTF�	B$�0k�"O4�8#�Ҡ/ �9E�.n��V�'=�����0t�l ��$^6�U��.>N6݇ȓ��[7G^]?2�Zq�j��,��G4��C^k�؝��D�f�����V���F�,f`#�,��8e�ȓ =Fe���8N�hH`��!@6)��&ܝ�FD:z(\�Y��L�'\��Zs�i`��<.�4��/���@�ȓ%�x4Yd 	2t 93i�8t	�Ȇ���mq&�2ZF�x�o2~���ȓ&� :�����z�8��-N�؜�ȓ7xx {g,�yhL=��/M*������2�O.$��B<Qi�s�������)&"O4����C�@��`����tɳ�"O����
s>e O�x|�ya�"O�Űqf��<��챱�R25o��"Or�ar�Ch~&�$�S�#YP=hA"O���6�ՊG�8�Q�F88S�����I-^@F�~Zf��cz��/��9(%Q%T�<c�^�L�<X�Ĉ�ez���N�h�<i�Y2*/4���r���xLd�<� ���ק5u.��OQ+���"O$�s�*�;���V D~:�9�"ODy��
�r�u/RVJ�c�'.�,Q���S�c���v�@$J��{����~}�ȓx����Ձ]>	�<�����FZ,���%�y:�e��Qʈ�����~ٸ��3��Y�2^9���٠4��,�ȓ`� 3�P�Cf�K�P��u��mu�5��Ъ��X�\��!�')�aQ�8��D����L(��!_=+t,������A�>1[�Lڕ�ٺU�z��ȓD�2�` ,�:fy��z���@i�a�ȓGΠxj�d�6Wcp= BO�,jڮ���L�6�
�K�1��Q������;n�B���sf�;�l�f<!I�L@,�B�	83�xR!a߽_��B�b�Li�B�I�?b�P�g�G!��� �?�nB�I3�z���ɯ	9��S�$9�LB�I�*�Vi #[���H�Ơ�1B�I�2"��(��C%΅z�'�f���=��
\s�OV�s���>�@�R���y��h)�'���7��"a�� ;�q���'[��� ss�a��h٪�R1p�'z�iG3^�ŨaIզ
�V!s�'��Mɰ��)�hy�E�x���'� AWi��=r���U�ڈ��j�Fx��	ܣ1ѶU��$� ذ���T �B�	qؘ<k��N-L�
�1��R��B�	 ]�* qDSq� �W�_�Y��B�I�ش���V�w�(��G���7  B��.L�F�P��OW�̔i�L=pKB�	)=0�1�@�d�r���6�<��=�`Ir���u>��O�$;�ε�CC��p��Ls�"�?"O�J��' ʥY�'9��'�n	8�Dсe�j�CĤ�$2g� +v(�º�Ѭ͒t"�� W�ؐt,�ɉ��Xx�'nDea�I4(�
�Q�;4�BEu��	C൩r��%ZƔ�m%������ٟ�|��̉#� �Z�o�>H��Ly��'�Ĭ�2��!h��(����۶� 	�a$��("i�dʉ����H�@J@ʓX�F<*���?������ʋ-����O��Q&+8.�jq��-N�����O����ߵ!G\@�#D�_HtX������i�7o����Nf7��j8��A�5p6�`���c�0�vÁ/Ywb��; ;R	L~�d�8��x��� m����M��<فIK��(��z~J~��O}�0��Z�q@.͎}��� �"O�ڣ��Ve�qd,ڙ� (����>)��i>��"E�X���(#$_6;nVm1���,��ٟ<)d^�0�.��Iȟ0��ןtYw���@1j<��8T$yK�����;�Ь���S�zF��DB܁��#��?��?)C��aB<����� LS$<���
<ZrAt�"W<X���C�<��O��O�� ��!',>0H3�! �d�"4��<�� �����ٴ��2=�H��c��	T��bM��Q���"`"O���E(468 ��4L�{���7�'{\"=!�i9rZ�h���ܠ}~u;(�%pEz�L�neH�Q���蟈�I5�u��'"<���ǫQ���P��bT��x��I�|��E�֭S�]"�J�Hx�����'s~I��e�76y�����_�ň`�� �vx�`��Oh0���� /�0���>^D�J���OJ�=1���
	#���I� �4K�!U8�!�7pU4\2a_;T�4Y���"f�I��M���d8j��OG�7�<{3Ճvd$T�A�;W���Rq�'�9W�'t��'W���`���c�ԛ�� G�Q[r�M�;��Y�޽+����;<|\�抗]�'����m�3@cx	Y��M��u���nݱ�ǈ�,�	��Ƒp����MH⦩����� ��ḩP���&���b�D�B��4���'�a~�lP:�m��&9�, �ea���>Q�^�<,� 1�@�:g�I(�ɗ*��˓M������?�����iA3���O0hd]�P�=i�ɿ^xd$&�O�us6���@d���H9ZI8�b������Iɴ�ăB��=4�0���R� ��$�'���Ѳ;����jE/3��|���u�E!���I�4���-p&���3�؋c���C?�������D��� ��2&��aB�C��4$ƚ8:�"O"s�Ϝ8RX�$!I�H\�f�I�ȟ�A����/(Op�j�ϛ�"�R�(�O����OD�q$�w�����O��D�O��;�?�S�3PNhk ��3�dA�g9쥺�+6͜aHp�<K�p!�˟B�0����n���cS@����;xj =�s�
�KK�E`G�Ԉ^T�'��'a�,�@�R�V�;�ML�+d��c�O桊g�'��'�O��SPy�(26���˅lT�߰C�h}�P!eD�$��Ӎ>f4�d�r�����'1�'�6(�E"������@E��
LJ���?JK�9��̟�������ǟ����|�A�hJ��i׎;I��ui g�4�~9BЧ��E�4e���6�0 �		.���M��Q� ��8y(8���K�)��L< �	���B��MK�4r~�OP��҅��	8d�$�뇭P&�<8���hO�">���L�H��YC&��;a�	Y��X{�<Y� 
9
X�L����Y������uy®`����<a�,���?���?�O��)��e�[��ś��O>O�:�k��`���?���� ��E�͍n�0Q�E�¥�?��O��
qcQ`�̡`!$�!	r�c���Y8gD.`K� CH�q�M5EB���@�<L�|�CIO�3�q��n{���'�O��$�O���o>���dZ"�!���*�ٱL�O����O���O��'��'��32lQ�?� ��fʓ?��a[��'�^6��ݦC�0'�&�pG鐼>8.��U�A|y��'��6M�O�b>�D�O���-@�H&���!)� �S|H��I:a"��{B��(5�,�{e��Aq�p�$��3�V⟬m�J�I�8w�O�,�p� ��:�I� $������p�ǺI���I�Ur���O�)�O,�ɾ�% G���hC����	SH��Ed�����	>S�i�I�<9w��tnz�E8Οk쒐A�:�:@�IkZP�SBG� ~4&���?������y������O��)�O��	�S>s���4)��҅g�H~ye �O���\�_a��p�C�	�?7��,�c�n|x�l�$ެҤ�U� ��a���5ʆ��	��2o�����O�����6��Û+�#�͓5t0`�%C��^���I;f�����ONȨ��O��ɴp��s���Ǻ[�i�3(G��
U��$!YIp��ڦ	̓]�����YD8���?��� �`3�m�@����1mZ<��v`G��y2 H��?��r��O牣yƶ�s�Nt�G�48��,ˠ@�H����~eĈlZ�<	�(��M��i`L���1O���?}�S3.Y��)˶YbL)�sB$u�|�(�4
�"�Ҟ'w�D����?	�'�?Y�'�b��O�F�jC��[2�,r�#�R�;a�iXA�W�'��|��L���݊�'��	����EX�+=�Yɀ@ҳ]~p]3���l�<��*�s���7��uA�9/Q�7��Ot˓�?�\?�'��5@��·l�8L���u��`��	Rڴ�?����<ُ�	��*��|��A#�(�AA�Z1+D�OX�O��<yE09�h���69I$4rtHO�<ACP1u1
�h`.ĳ_0����M�<���[��	��3x!͙b@�G�<9E�B�1 ��q�h5}3�M���E�<��W�rZ `OX%�h�n�Y�<��E7Y�<h ➅"�E(B(FT�<Q�l�l�`|��F�:琝���w�<�F yD����G9�li��I�<�P�ؚ^���͈{��PQ�m��<���͆0�vU�e�C�7�����D�U�<����3q���������1X��
Q�<y���f�F�1�k�{�����h�Ak�JW�t:��0&�4��* ݟ7�L�gB�zy�6�/c��D'�nцa�V��f�f��L%C`z����;V!������S� �R�V��ՃΞ&��|�%���N�K�i%+�(
�m˂W6� �pi��^d!Q��	�^��D@�1�%���dJ�>^�d"��N~BZ�%�!o�!�$ݴcX�����?|l���Q�	�!�V=f	�:��Ċ�����ԹT!򄙆ԺH��M�}�Ҕs�C�s%!�<Ҥ�B@�V�4,;7&H�!!�$ڐΠ�Y��
�%�&��De�w�!���y�x��㟕�f��p��<�!�D��)g@9�U��E���2e^�K�!��ƀ7p�2`gN�*���j��ڌN�!�([��dk��~�T�x#.%g�!��	��3Ј�$�� s�mԑ*�!�D@?��k6O�N]=�M�0�!��i N��5��)��e��W�3�!�� (�25ʗ> �!�d]0h��X��"Ov�{�hP$�$�TNߠ� ��3"O��ip��&]2��׍� �qҤ"O���e�D!`�d���*F3$���:"OvX0c�7� I�i>g��PHu"O�Iɐ��2#~F0�$�1p�*H��"O�Ճ�)#���aFE.q��"O��4�Ca����#N�1�T-X�"OZ)���)S1V	a��0^FX�"OT�� ��0K�>���B��aA\�"O��ST�G���o֩u@<��A"O�� 5�@��e1@�*	.nPH "O3g��|���5�*.+|ɀ�"OR�x1�K�D庄�2⍿@���1�"O��ꂡ����Ӗ���pu�"O�a��Q!
�T�%��}�ް[p"O.����2��T)�@Ƥp�x<8�"O�L�%�)��i#�Wk���d"OP�� +��b����웘A�2�K"O�YE��p�P�y �#�f�Á"O�	�d��0
���7�µ!����"OV���:-�ݻ�-��1�f�i�"O���E�	�x吃g�0��)X�"O���H�����r���-����"O���ɒb��b'鑂S.��g"O*�*o�1�����hN�/,�[�"O
a
E��:
�����8Qȡ"Or�H���>jRP1�$͔��e"O��k�!�� f!���\�����"O�	B��ʸX�r��(����I�"O�(��U%bn"lH'0��Qx�"O�,�&�q������P_̐�"O
\8��&U�w�ˡS��q"O�p��Ҡ!��(�+PP��]��"O�]1��]N��Ҩ]�8��Љ�"O �AA.T/�N�9c'	� YZ�"Oʍ�&���(��	1�)2?t��"O.E����*�6��B�JG�q"OX��D珮,Ȍ��SC�8E*,���"O�"�"�k|X�[�`��S�-*�"O`-I��w�VŰ��i��+b"OB ��L$�E!�.�'5�b�k1"O�}ە$G'}
�+�ML�0��(��"O\�3.�sv���V�j)z�E�<a�hW�#���it�L��(@�&��@�<�Q�I�n�"���4ސ�`CQ�<	�dA[
Z����A@I��i�<1A�AE�t���-Zu$Y��� O�<�L�)���(q�ߗ5l0(�tH�M�<90�7Y��� �nR,�@�bτT�<5�H*�9" &�%Qa �p�)5T��k�Ɯ&&�Z�2��c�q!��7D�4�W�Θq`�u F��_����1'9D��A��>��ıW�A2@��$�Ѣ4D�<Z�f�,�e �c�(�$eF?D�Xc����bϊ���NT4L�����=D� Yr��d|d����R�X��b�;D�H�p%�6QB��c�b�P#��:D���3��	�hAP�

�/@�]��j$D�<�� 	��lS�e�+'�ᆃ"D��5�g�9�tmE�I��ŀ��$D��#EСL.���%A��VD�ec$D��Á�]�����`��%l�R��G#D�X�U�� �!kU�� (pW�?D�� �ժ5�P�e)LԠCCуj�(Z�"O� �d��v�Er�aO{&4� �"O�9�%�]
D��9�c` �%�"O��tΗA3��x!߾s>:�۵"Op�#bԫB� �s �D�1"O��`�r�!�.Jq��"O����`��@����D���1A"O����ɒF�
1��A� urw"OB�Y����BXU0#%�:ax~"O�l� �^��Y�TJ�Np���"O�%PCh\bbL��=m2���"OBIF�bl��v��/1c�"O�ئ���h�X�c���:g��P�"O�%��9mĮ���'�9Q8�2"O.ũCI1S���Rȃ�8NT�Y�"O�E����;�n��uG�*0dT�"O�j��R���l@�F=07\�"O����L]}������:� L(�"O�JRn]�B��(&�Bˮ��q"O�=ѥnZ�aUZC��0QB�"O4(pd/��S�hR��p���"O�آ��	��A�ڑt� M��"O�����%p����Dj��&�*�p"O�ݺ&nQ2g�r [�iPm���s"Oʍ���1B��+�ȓ�>���"O�\C��Y�L��5����D+���"Od��A�r^��&�v��"OȔ@fO)c#�H���"I6<b�"O���!
3Z(`���GHjpv"O�����8C^���/KZ+Z؉U"Oj�j©�Fк�� /Ӽ�I�G"O�`�a6D�)S@/P/]��\"�"O��Jb˗5�t�[��L�+� i�"O���,�Isj�3�B��3�H8�"Ol��kʛn��H��g.s2�"O^�@���	C��UZ$�Q�%��l�R"O�Ԑ��n�zг�F�\�	Ѥ"O^���>@+<HH��ӦP�� '"O�,s�"v\���jRv�H ٓ"OȨ�\��*��t�!3��B!�dK�!-J���&M�p|1��V�O!�d�l԰q�GZ,�D�d��b�!�%Y+ )9�� y��T)�뜎S�!��ɏ^�蹑/G�!����!��H.T��2g2e�t葤�!�dS��@�G���ݰpJG$�!�$�H�,����r�<�F$��yg!�1a�5�R��}�|;��F�%f!� 
�>�SŔCf�(z�#��E8!�D�'J�,T�Vg\y�&�0�d�'�!�Y0IS�iY�e��r�� )qɐ �!��R'2�V��� m�$ٓP/�#z!���m.������Q�e.�p�!��>>=RpZ���U\�큳��V�!�FzDɦ��@���uMP�#u!�$��c� a`����5+���Q�;GW!�D��~5���'�(&���]l!�$�u��A�.1W�!Ӱ$H3d!��Q�,3�eA��% �PA��ɣ@Y!�$���^y�g�4 f�j%�	'!�$"�v��'�V�P�L��ā�,�!�d�D[dSfO5C��0�d��u�!�d��_�������qϮZl!�#˨�YU
�<���S�ҁZ_!�� b�r',�>�xD�*
�X�"O��K�BЇ�"1�䗍j
���"O�ab�?�������R�U�""O�a�G,�3D�v�[S���^�[""O�1�����.Q �n(b%Pp�6"O&�1��-�j��+y�e*�"O@�y!�
�r��+W�E�)��"O��zP)��ANP!�!�	Pf`"O���e`_2&[���� �;b�4�9d"Of<&��
@	��ڹhL%�!"OL��T'ؑa`
����_1d=0A"Of;�Kb!���7G�Е;TBF9fO!�ą<�X�dě%aN��S�@RM!�T.W�#�ϋ�P<,���E�z(!�$L:.���"p.�n����V�>!��J.tv9� E�Uc\��7�ދ4!�DB��P�`Bȡ#3�l��S�!�V 7:�������Dz43���	�!򤇯����7-��!7V�r����!�d޻$ I��fK�s.r4#�(�	j�!�#[>��"qBVW�ĵs�4a�!��ן�>Xa"J�m�H�ȕ�6cC!�DwJ��f��5y�*��2L%7=!�OPA�$�%�L��aTJ'!��A	K�(��q��4Cɸ�!rbν"$!�D��i�z呃4���)FH�\�!���(�@pca���sΔ'I�!�K�U� �H��W�G�|\��sG!�D��]��tD4��-"C��2!��G�v��t�чʤh��)�v�`!�=0=(���'�.4y��^�!�dB���a�e�^�9�XH;��ܼ!���8�8�i�2�i�i�'!��9b#�A*� �t�ۯ3�!�dV7+	Jzw��:�����j�!�� H�v )S��-#0y�eǈ�`�!��Z%qk�H�Q�A��BS��)4�!�(0��qQQ!�8<T�  �B�!��̈PY\�[���%1�r���1 o!�$�X83 �2a��9KO�!�$��}ب� �"Ż>j���J
 G!�d +t����%`Jy$��KS�^0!�d��>̮(1�D�e� �
�"�"~�!�$���kB.ɮs����e�� !!��W�x������Lj����3�&�!���0!�\1q�D!�P`�O�6�!�d�=t���ҕ�\�@�'�!�$�;UƜA0�N8}�������� �!򄗤���X�f�!��A��!�$X0b�B�7&��3
�����O�!��+�$P&C$V�е�ݤ�!�dٱ}�p��M^v%����='�!��܆x06��	فZ+��d���E!��N�~xɂ�ĳ\���P�c��j�!�d�6�5HĄ�E�1��+�!��"�:�څ�O2|�!9� 	'�!����9��`G  ��b�,���qOʰsB��0��$q�Y5&{J ��G�m	�X�P��9h�%ۏW������y��y��'{�{�k�6�N$1�HlǶ%ʱ;�l!L�lI��<Q�"��S��R۳4�N=kS�Vg�<!��$�a�fG��g�>U�2	�?b.̠C��(�䘆�IqJ�*�L�M��A�HŪu֤��dC�7P�P�b�U?I��ř���SH�B��teQ�<	�□;��qɵMɝLO�3'.
oܓg�G�U7Q?� D�2hH�;���÷lM�m@��""O�kw�B3������L�0�����6 Q$����<��ɧV"~y�p�IȬ�ӒN�M�<�DH����,��l@[�<|k�/�L�	z�Na}¤,!޹�w�õR�r}�v�1�p=�t�ě���2�m��.[*���a`��&$���t
�qs	�s�ļ����&/�>��=I�e��#j�𩊖$�y� aH >�1xT(�j�!�$س#�J��r�O1%��(��J�<�?�R2�gy���8���ʑ��t�$�Sf���y�E5����+��d�<
�[�wq^U�'��B�R>-\:ia��[�k\�S�'��X���=wk��p3�_�Ԑ���U�oȏ5C��c��X�n���D�-D�\��MB�e������b�8:�,+D��� �uc� H�Ł�d=�#+D�0Is�T�7�|�#E�b4D�aG5D��K�G�B8, 0akƏnr�%��n D��Ȳ�6�YP4�s�����-D�p�L^�2�d�����9H���ї�/D����`� ���$9'q��S�h.D���O�.3�
P��?x�f�T�*D�hy3�]<&���4���#��x��.D�l��~�K��֮�<`yA�+D�D�B��[����F֩�I�po6D�L����Xl�����'��Q�3D��1@d[���N��]& %D�@*r@B�5�M�	 �V(��5D��2���(%�e��ݵ?�\��7�(D��(��y�򁙦�\"�0%�F 6D���'`�5Cʦ��Q�\�T��Aa�1D��j��ي+��ts�K\�E��pw+<D�<����#( >�I��E��0<ʓ��<��: �|�+���jt�
%Ah�<!ǆMJe*���I�j3G�Te�<�`�&66n��T�
�kol�(��b�<A�'�v�L��H�"5� ���{�<)ǅP�A2�ic���O����)Nz�<9���)7�����֡�KL{�<��4�\�����2?h ��n'D��aR#]�4���ҕ���I����U�%D���$��'�����)�0kX�Y5�0D�t���؝.ېu����K��T�$D���p��W|>e)@���0`�"D����c����V$�T���B� D�����*�ȒK� ��dSo!D��P����_����_�!X�UP�M$D�<(�"�}�8Xc�g�p[�iF�=D�8��B����4'L&f���%c>D���ΐ7q\� ����	���yh)D�$���I0_8<T�N�/7`�a`�5D����C�>^�%��AP.Z b�hF�'D�X"`�U�
�ڤ�ߝ���(0D�H�w�9x�89��b�#'����<D���UG
�/�&���	sw�Cn<D�p���5q����΋+JY��Q�o8D��P����H�ࡍ�u�iA�d<D����G�_��-8d	�%qT�z�!;D��i�Kܠ'<J�+&C�;��Q�"",D��	�!
�%:8�aĘ" � ��j/D����H�5���f�L���#-D�l���3u�$Ђv*�;,JT�%�(D�ȂF	2|A��b2��{O�HU#D��q$F �xУ�$�'sr�}9')!D�� P��a�������!�k�\��"O�ă�&�1$Hz�'W6�1ks"OVX@���9O������]b7�Q�<	���w�k1?GE�X���G�<'D²!��4�ţ(~T���H~�<9��^'N��t��ϊ)$��1rA~�<9(U-;�"��'� �*QD
`�<� ÍJt��yq)�r����g�Q�<!`e̒{X�Qk�e�r���Ӧ�C�<�����9E�jb��&�
�sP��h�<y���/�b���Ɖ���2M�g�<a#�3i?Э�FKEE� =!#ICh�<ǽ(�TE��ɞ	�ɂfQe�<�f� �z�W��)ݨ�Sr*e�<)w[`P0kF�7J�j1��H�<1]����7Z`�i�uK�I�)��R�!�l��WK��
V��*��ȓz8�1A���,\���
�-'�U�ȓW=��'��(]�"�X�LJ-�ȓSf!��O�D���[%Oـ>�ʁ�ȓ2�Ԑ��fn���suA�Q�|؅�4xx�`DqH)�&n�.�>9��q~��'�Q��M+�f((����D�X��ʊC;��6b	�����ȓ<��y !c��a�b[�{�"̈́ȓ/pm��V	m*�{T�J�w�.���r������7o���S�H�,B�L��yvހ��'ْzԁå��(��ȓ8�d�8��OLr놃	�E�1�ȓNE��5�����|(vmL�=���$��!��8*/N}�p�E��V��u�R���̌�E�ʑ���S�u�D��ȓ'��@�f�>�F(ҐDB��������*�bЏ"�xUѵ���r�
��ȓ!=X��AGP�0W���ڕ]����V��@��R�t9��hʚ	��KO�1����N� :�j�? �P��ȓW&@�A�iΨ�kT�g�&���u�0љ�]�b5��A_+B���,kn}k0EW�@Zl`��Ly\��b�������eB-R'ō�(���ȓu)0=��|X����� �,[�ۃ;�JH���/�m�����'ej�2��$�dlj���51�n4��'B���cB�[�&��B>��ش5��LIqo�$Y�h�``�ϯR��G~��Hfmr.�3l�$ɒ�	���0=	���X��IˀO�0E��T%���Y��KE��L��E�ab����'�|呴�E�y��(:B��nk��P�yB��N+��Rq�G>	�\������M'>]�KA��D���A,����=D��u�tp���B
�z���#s��@�D�]��a��lcӮ�G����>9��ɥf�D<[�l�-_����qn�@�<���6��l*��߭��,�4�A�� �nϰ%������EF<j#
3�A�Є��'f��0�"]�2f�\��8@z��C9sʮ���Um�d|q-Z.c���pT�\�!����A���?YqJX�\��`��8�"�l̓�  ��U'���!)�.HV�Q�g������� ¥v�@0*bɑ�yR�۪1��d�$�ٽd4l�S ß9����]
B��IB�VE������	�o}"+
T#��bP���h@s㪊��y2`��U0����HS
����ȦK�v�[�X�~��U3����/�m�0d'�xi�uI�.��3�<����
4�(���	p�ti��a:F��I���.o~��҂��t"4��Ń�#@�H���oK�?yG�� 3���y@��<�P@V��b̓�PAT�Ͳ7��0��ٻG�N��7��$�E+Dנ� �O��Ohh��)]�y�T."��Y����_���#ᎆ6n��#6D�U:-��ax�nii��I�M}bć��eȃ�֯]2�0��$�y
� ��S� �z�I��/,nq �-�5L�p��N�D�~����']�F~��мN�\�*:G�p�@%`״�0=I��D8|��cJ|�tH��0�`��!�;	�J���k��tz����'7��AG^�*]s���/a~���y���!���pKK>D���ը�0�T����P�L)�H<(I0�c"O��1s�sr��-K�T�<��
���9C5/(?Q��K��i��#|�S���p�#�d�K��t��
'D���T�P#|�&�˷A$8��킥os�jk���$:y6�� ���0�l����� ��A�Oyc=�Ќ�V1B0���61̞|iDL�X��
��Δ=:X��,�8�akD�Z.�6M۷��5��?�HQ�����)�0V�l�०b�v���᧢h ����=�n:���e�p�NZ^(��P����N�!�$I6=h|+T�H2 ����ӥ<�d��֗��"'B�*雖�;�'o��� Q!d���N�UÊ`�g"��C��+u���[&吝y5��vDX%��6�V�$�1�@ʠ ԏw�����W� A��S̗<����%D� �EGA�&�(q� �ٴa�vt�+6D�0�E�h�hh��̅0%�̠�� D���f��xe�I��D@R��y�(-D�����2�F�͑1\�;E�*D�������dA#Q$"d�����.D��(Gi_�v}fe���6J$�|��B-D��HӡA�m�Z�f��S��<�9D��t#�,]?�=j�M����*D�$��l��S���E�!�*D���Z.ł9�3��v����2�)D����X���e�F��|����5D��H��(X��3�X$�Z����4D�S�I�>I���������,%#�-=D�����N�"hV�]�Q�a�'D� ʀ��|4@�E⓸h&�q+��%D�d[�n4z��T�2���;��y@��#D�$!oN�>�>l�������z'g#D���#遆���LՎZ��$�$N5D���6jZ5V.P)�I�H�l�K��0D�������)3�Q�j~8l8# #D��٤{�)°��y��(�!#D��viEA
��]|�z4���!D�x�����p�K"&��.�R�%D����Ğ3F�4u�6O%R��ը��?D��У�f�\�R&�}E�0��=D��a��Ϥ�0So�sy�U�֤=D�`�o�89Fr�@�$��ܝ)R�9D��@M�8!��yِ�ա7�� �h;D�D*�jH�kl�mA�LӜ%p8�� $D���a���a�b��2�_$`9�}zp�7D����ŀ�5 Hr��\�=Tqi�%6D��S�O
W-<���l�%pN����6D�x*F3~@���VÛ"I�:t�*6D�4@ZQ��c����b4D�Pq1��x�Hg��(B������0D����'Z@�zBD�LMؕ�2D��K��3:U,���+�h�j���%D��bDҶ݆�27��7X�B�J3�-D���fe�7N��m1��ɆF�b*D�0v�� M~`p��̾Z\�M��)D���D�I0��H{E+L8lQ~�i��,D�ܨ%�g쀽`2��RH(I	�,D�Iv�
:E����-�3�-���?D��SF�Q���Kǋ��;Ԟ�!'"D�H��N�<>vԩ�!I
��؈&A/�	�D-�D��C��VZd�Ji*ВO�T+WiD��a�@�hJX�`"O��Q�@�C��д�Q�	��Z0"OV4A�!�*���g�!Y��QBR"O� �$��Ʌ�7B��`B��n����"Op	�r�V(��}`�hZ!H~�T�"O�a&@Q�sND�c��ޠkpX�Bp"O�P��"�_x��vힲ2Z��A"O�d�ħ��,Y���I�`G�%Ja"OPeRaH�twJ1{b
*k3H��"O@u۰�J�4�dm1uIT�(8���A"Oօrc�Q�������:+�ܑ1"Ov�:v䄳!h(�G͂26�@�"O�iX 	M"B�l��+IVp�:%"O0Q{1+�4`M�܂3�MRAҥ"O@�{`�gc�Ҁσ���:�"O�lcM��l��в�����!�"O>xx���hiur3IӋ\E���"OP�{�A�-d�� 」�R�:U"OB����͞������6�P�Ba"O�l��e�������0X�$��c"O\�(S��Z�|9*EL�3xzڄ"OIk�H��8����ǲt[���g"O�������^I�	�#�W77R�С"O`���H�.��UC�F2�(�"O�B�e�Ju�U#F.k�"O��`�H~l��XGp�)t"ObAf�H; 3�ɀGX��^!��"O@H����:p�%iE� ~�~���"OP��E�6�3�!��$(@"O�DaP#B 5<4{�m�Q�`H"O0\��\W�������$=�"O蛲�[m�>�"	�0���"O��a��jG���`.���Q㎯�y����{��E� CTT���Z�y"�521f���ϟr� ��RM��yR`��Y�\Jefمc�Z8Rc�ւ�y��U�L����4L�h�&̃R�y҃��Ty�q�ġ	=����Q	ľ��'�ў���T���R'n�b򡂍k{ʌ��"O���τ!G�ZF��t�ʥ�B�Fx�$3�����RUI�>h3>P��-!D�Y�ąkn^E)���:Z�eq+;D���%�ŨQI�)�H�&?��6D� ے
I	�	I�oմn�d�Q#�/D� Q �����Ҁ(A�,B´'.D�H��#�0*uH�+���x�&@ygM+D���+@E��B�]�k�*D��{�Ʒ$	۰
�&.��G'&D�`
�!��ݖ�9�.^
F��x)�('D�\�dNݱV� ȪL�M�0=
�&D�D�e/��E)E�G�d[�3��%D�cTH�'����q c`"	q`�"D�H���nJFtRC�#,`(у/;D���8S���'��q��[�C9D��wK�zV,��JW%2���6�6D����
L�|=t����G�&���k�<S�� z��-�f�Kw,(�(tf~�<1#%Y�4|6� ��K&Q8w��A�<a`@2h�iS�bH�j]*I�C@t�<�5��#���Ԯ��z����s�<y�#�Cc���ǒ �H�GaGd�<Yqk¦��a!�@���JSc�<9T�"��p)��rm�Y��]�<��nX�XC��6��0�(y�fC�n�<����8�h	�M@^�:��^j�<)!�@.ԨZ�⓭�^d�Ef�}�<1M����IB���|��8J7��|�<� n�ʖ"&�����ǆ�3�~���"O�)���A_$�p�ص:�ᐶ"O&xH-�	�E���

t1s�"O��c&C+���u�ڸe�y{U"O<���#L�c9B�
T���J�l�p�"O�L���=%0�a��)%�zɊ$"Oܕ�2��+~մXڥ(�b����d"Ov��	�$t|!3v�ͻ��Q��"OL-sɛ�rg>q�UH]�{��9: "Ob��a�^(8ՊF�1h����"O���с2+L�
��FPM`DS"O�����=�q�KL@Ӓ"ODq�T�R1�Te`���OI>�0"O��pm�U�8P�%"�6\�x7"O����,A�;�:����0pf�qh�"O0�z�e�Щ�φ�O�� b"O�kp�'w>h��W;;/�1qR"O����B�O_�ͣ��Yz�]b�"O�}����KHpy���ŧtg)j�"O*��1�A�-B�9�&
�	_�$x"O|���
�GD�4�`�+!�E�&"O�)�G�"@p# K�O�	�&"Oxm�BEPU H�I®��F58"O��f&�(���Ʋ"W�DrE"O�������7���8&%�qi�"OZ�U#@�C�X�[q
I�r�0i�%"O`p�a��+��s4����|db�"O�$��M-��I5��%@5z��0"OvT+�`�r�=���#o�Lj�"O�de]�,@q��=p����"O��S�g��HУ�l�f(aA"O�]*S$�/*P( c�H�l�b�"O�h�"�<6/�yу�'+�8�"O��!�k�y�eꦥ��Hyx
!"O�93�EP}���*'�׼Mwa��"O�1G�D!dX�%[� E"c�lC1"O(�U�]���ə�¢X�b��"O�M��M�;j�2V��bQX��'I6P.�ha�@٤!�F�8��]8�y�a��I<8�+�L:v�0eF�!�y�V2eT�ݹ��'(��0a��y�ӻ;���`�����`���y�J7v0�FNðP��L�y2!_��j�Ci4!�G����'�Vi �h�FǪݒ�kTx��'�2��l�6N.,�SrF�.>�q��'Ӟ4`���"ew"8�
ߓ7�����'9�k�(}V6�r���+����'��y�EA�|�xiT-X3 :�i��'��M�M�<k�fx:��W�A$5X�'��82�ߙ7R�S�	%��]��'��]Cp咱R���aQ<|�mB
�'�f��6	��T�0��@�7�P�c	�'ˢ �E��u���*�:z���'T���$P?P��M�(�+2@���'Dt�Ҵ�=��U"��'z$(K�'�`,Q'�?�����e��b�'EH����_���3�C9b�����'Q�	B�(�'H$f��B W����	�'�����I��!��`��>4:	�'��:��3q2��!��`���'�~!��ݖ/�"� �&D"*\|
�'n��V���?��}Kp�=\�LL�	�'3����� _�X�g�С=��9��� b=a1,Q?*��	�Q�V[j7"O܀���*�8w-tP.q�$"O��e��cc.��W�E;^��w"OJY
'J+i����i�hn��C"O����tF|�)��B�9�"O.m[ (@�$s�AS�g*7�8}kt"O����2|8ͱ�� c9�%{3"OD��bF�`��2 #��"O��h����YB�+�d�`�"O�%�1�L3u�a	����4���"O��0�F���Ik�
�]�(%��"O:��Uʁ�Q�����L_�H��ԡ�"O��i��6BI�J�k\�k�j��s"O�]H��^��4Mg@��r�옹r"O���T�H-��0 ������R"O��c��:�\A�jح�x�t"O9��6v@!@���Xp��"OhԂv����I�!�+~Y�}*V"O� �wkܭ'�vdcS'�i�.�iT"O��'�
�LyzP�և�<X�*Ո�"O����P�&=>�;�'�QL��7"Oz��J��?�E
���.,U�$�b"O���tТ�+W���{�|�W"O�E`��;���a/��o�n�`�"OFx �
�u\2���Ν�g�>��a"O���u
N�G��hquo����2�"O��ca�#+�4ẵgϓY��h@r"O�)��HQ!$�*�$�ݨ>�p,Á"O�h9'�-D��4	C�)	F �"O�@)pՊRN5�AD�:�F@3�"O��Q
F�/-Ҙ��"ܻ��X"O<�0����LT��9�����4j�"O��C3c7���'L�h�\4�$"O.�k����/;r��kF
�8��%"O�BDN	1�rD�% ��[�,�� "O��GM�g"�5�Bo��7�h割"O�b凋��`��ۣ(tPd�Q"O��!&:������8h�-��"On�j4"��[��hq�M��*^�k'"O�$��%Fjz	��%��\WȰI�"OR�h�O�f-h�n̋Asr|[�"OD9�#Դ��$��À�#�"O\�S�m�.ذӰŶ	��Z�"O2-A��Ɨu�\̸�+�
F��"O���Hb�m1�Zb�La�"O�IQ��^�/��4c�ղ��0�"O���W��|k� �|��B"Ov� ၀)X���mFd�h��#"O��〭�ry���C섋Z3^|�F"O�u0�o�q�`���I	:4�"O�Ԫ�jCX��đ�`�\� �"O�u�aџo��`r����8y���4"O�y{ĦVג2��-���`�n���y��О.�<���ޯ"�&���Jա�yRB��Q���&�#���# �+�y��Hp�c��
]���ai��y2n� \j4�����~w� a,M��yb�֣Ij�	�Q�3E�Dc�&ۛ�y"�ξ�q�'I��@�5*T��y�dOj=�L+B˜�4�9pW�	+�y.�@2���Ԡ�'%8<M��ޙ�y���4 �
&HH*�x�/ӿ�yb��JE�$R�O�x\!�'���y�Ȉ������Q�	�w��y
� ����ʢX�Yz��ʗ6�~ �V"O���3<<p�I�&��2"OV��
�6ED���n��Y"VQ�"O� 3T,�E�`�Pn�)>=��j�"O>�;�>���e��z�"O��sUaE�7d����Z%A���r�"O()S�˛�xN��P�dV���R"Oʱ��b�3�B�ڧ$zE�[1�X�<i��'H�b ���	%D�m�F�x�<16�
�e^ �� �m������M�<���V�^�6�{��3Q���l_�<9CC���)�����$�A�/�X�<!P!كR-�$�VE+w&9� KQ�<�҆�t���b�7y����$SJ�<q��$��Ի��L�n��P��@�q�<��I:���脌I�8����Bs�<��A�f�f�a폣*8e���
d�<��IS�	�f_ILP���J�<�4Γ�*b�f�W���'�]O�<! �At��t�n���T�
�`a�<91��.�ԥJ@͒o�����v�<�ԄS�������a�F�����i�<Y��I%  f�� m5^��(��c�<	�C�b}��㑊�.zd���]Z�<	� C�W!ir��X��	�Lp�<Yo8�Xx����d�zS(m�<���@�z� OΧ:=�`��+p�<i焝�{�d��'s�Ȩ��Q�<)���$)��9��HX�X��\���M�<�ǘ�)��0s�ᗗn�ʁ3U��o�<�
��{n���g��()��k��a�<Q&�$�X� �EC�-���y�<	��W*�<	@IPY��zV#�r�<��(M2Q��`b�ϋ�0��}���Sq�<12�H�De
4r��̎X�X�n�X�<��f�&1r��F�ss Ez�AQ�<Q֤�7<Rd �l¬$� �١c�L�<aVOY[����QD�~�Y�Dd�<�A��I�]�wW�w�RM�"�E�<q���!Az�(�'@Ŗ Q��@�<�5��!"�E���Zd4�Xd�F�<q�BN>�v\�Q9</���IE�<�u��;]���"��m*\ꅣ
A�<�bg�\d�AV"x)*@���$-�B䉰01 �ꑄֻ'k�@&dP�$x�B�ɅB��U@�H�".1Ѩ�М[�$B�I!P�\+bj��<�t��܎b�C�I c���H�	!�h�����B�I�c�~Q���J�I���P���J�vB��t[�1�!*B�����E)H8EEfB䉊����͏w*@���I��.B�	�_���R��rRa*�HB�U���H��-x�k@%H� ��C�	�6����!J��*kFnz�C�	�lq �W�B3jq:#˦Mw�C䉞Kv���a��W�d�I�
�f�"C��#�Dj��9�BM�`/J�t�bC�=�n5�4�=m��*Ӏ��4C�	�Uyjd�*�zs+-�/);� ��'&�T��K�`P��#��)&�*%8�'�L��Μ�j��t�"T�U%|��'��X���S5���_�`�fi@�'u>�01��6:�t( ����V�����'�8�� �#�T�R��Q�6؈��� ��� �5�,��c����"OtS%��|�J���K()nƩ�c"O���
L��J�S�EhhI�g"O�iBO	!S�pY�i]C��@p�"O� �MܖXh�E�F��o��@{W"O�Y:�&J%5��G�֥��"OV̠��B=W�XXx�!�n����"OpX��k��T�ЀS  �~�=8�"O�u�&끫g��L�s�J�2`�<�3"Oj�c�'X2J�x�n9b{��S�"O��x`��4��	�uHT�%]�"Oڭ�f��E�>M2�g��;MH��"O�蓤F��R�r�Ë���w"O��"���Kj�4���֟�X՘�"OVy3A�0)��&����1"O��㧂U[rvPQ��b=R�w"O���V$^5�>�������p0�"Ohj EZ1Bծ� Te�9}���R"O�ժ�� �AS���w����"OT���뉪z���a$�l��"O��"�gЭo��k樠���`�<i�&�=[`Z�j�E
�����%X\�<yQ�@����P!� DEk��Nc�<ITm�) �����ÉU�p� (d�<��G 4�,Cr����ʸ���[_�<q���g?�]�b��E�N`ӫ�X�<ee�5&��pRiO�[8 `�W��Q�<�w���'6��{Ɖ�/-~Jl��f�E�<��HՄ>@dzs��#0��l`1��z�<�b���B�]�Q���"�C�E�l�<Q�&K;h��=����?[>�ڇ�e�<�tE�5:���z2 Z�
�%_d�<ٔ�Q�Ș��E�K����	Y�<A�`��sܞ����~�Еаe�O�<��"לr�L���YK"��á�f�<q�������fT���UK�<1��r �jq��W�JI�S�<�$���1��#
�f$���wne�<���Q&��S�J�r��˵�Ga�<���K(S����&"���*�h�<	�+6)�\r���9.��q� �`�<atgĐ*��S�[�5�PqƧ�Y�<����>zĨdi+�0K�@ܐ�ǉX�<is"[�q�$y��
�'��e�,Jj�<�TgҼ��1"u��Fy��Ѥ�	L�<Y뉚eq��[���a�f���F�l�<�a���Y����G�#��I����f�<9у{R�Z�쉨�`� �b�<I���?��3����wX�}{�VU�<�q��1km~����͠v�R��j�<1�g�Ά����V�3���CnMh�<�4Ś%h��B�؍`�҉�B�BL�<)"�%/N�y����1~�x;$�J�<y k)V�{��۬x�8����C�<A�ʜ�u �$r��-^ƅ��H�}�<��ǖ�I������P.V�!gh}�<a�釫.����Q��v��Ǚr�<A�`P�n�.pـ��`_H�3�� J�<y�Nӎz�9�?|�A�U!�k�<��-H"M6YҒ��.{`���l�d�<��ȉ�L%x0�X8Oc�h10΀X�<��ն.@P����W)t0YD�X�<�fФ?(n�d��"��t�R|�<y���51��%�P�z��(z7�[M�<� r�7l�=bB�u��(]�W4ċ1"O\����S�"���0�JBvb4R"OёP�����i�f��<�z��W"O�%��JB4����?X좩�"O�y�F&e����T&M�~���R"OJ�e��"-�lp����|u�"Or)���F`�P��@�J�qm*��W"O�e֍_:[ת���ӆQ^`d
P"O��%�J7!�\ �bi)Jf8�"O
����g$N���I\�+K
H��"O>YS��޻�\jr�L<�Ƀ0"O�]Ief]u�3&�p9)��"O8�Ԩߍ15�`�d�<LZU�C"O x�6MN�Di$Zb�C�I��"O���S��!GgH,�U�9�Ƞ��"O�D��H�?�����	\�_�Lh�&"O �k�^�ZR$Sh�����p"O�3��4e�@�Q�W/?��M8w"O� @�
J�v*7+R�6p�Cv"O>��,X�mj��J�P��E"O(�+�8:C��֑D;T���"Oʩ惆dx�#ԃU3)<��"OPJ4�� ;c4#�	' ؼa��"O 5���
)�EZ�Ȱb"O���a�31ʤi�V#E�+��B"O��RN0{'��r@��:I�g"O�l�%�G^$��ׄO"
:@3#"OU�ir37 +�tX��"Oh=���Hv�Ry�BO�K���"O�1���_!�١d��t�Q"O:t�6��&0�1��61�Ω�g"O��'�0�&�K��#�X�)�"O���.�9����f��#M4�˔"OdM�r��n������?E:$	�"O���R�^�[Xj '�/U1�ɦ"O��3���MwT�K0F��/.���"O()��O
1BTt�"'?^�|T*�"Od�#S�&=����:��`�V"Ot�G��=,��!�D�;8����"Ol�#ӂ�	f'E;@cº2����"O������|�,�Pga��1��(#"O	Y#OX�[д�W�G%����"OD��3�R��k��˔�h�"OPd�/+r�a��%[� �$a��"O��JU�RÂ���đ�s:"t�G"O~�ٲ#�$E�Z�K���d,�He"O�x��.(����f���@5"O���S`13vL5�3hHOm�Q��"Op�b�  ��C,CX�p�y�"O�xA�!_���KCB�%�T�I�"O�BՌ:lM��[R#�!��SV"O"�ʰ��xs�kE��)v^̹�"OސЁ,R���	T�]pw�b�"O I����ooN�����kj䅒q"O���/ƣ=���CQ+\4���"O`�(�M.X�>�Kʆ�ò���y(ڟ��1��b�1��$�*�y�B�;�<�Ic��	�Jq�E��yR�S�"���6z��2�b���y2���P�yQ���=������y�̕�t��T[���.׾t�����yr��!K���@2*�,o����͓�y��	:�����?t4�� Й�y���
n=N�{��+ Qbq���3�y
� T�j2
�
 �̒��ɂ<_2-5"O쐓�Ɗ��$A�M�-#�A�e"Ov�QL
9QB`��t�+��т"O���f��W�eq#m��mi�X��"Oೀ�5l��#BL�" �e1��� ���^�hЛ��'6��W?9A�>I�*�*�A�UB�Q��.�k������?Q������I�z�j�� j�R%�c�z>�Q/\iR���ʅ(�	���:�O���t�����1 �� �J�+��O��D1fC�~�:�	���!n�@�	�%�M�'úĀ��?���i�W?����<)���a����8My�)��?�����'9�毒]5��Br�Dl�Ɏ{��	��M�6�iJ�f�Y�B��Z!U�� 1�~�j�����'�"]>�y���d��릩
��Ñ'��D�_+W����Qm�*(9Ȉxr�H�V6��[VM�,��x�qA�?	�O7��Ƃ<����z���bp��=rh����iVQ-c昘D� 'wQ4�0�+6�^1���\c��@:td����D����4=w�T��4I��l��%�MӦ�ip2�s�N��&�F�8�8�P �.J4`	��Oj�Ĥ<�
˓k0;u��&-��0	I�j4��Gz�i�6� �D�~2�f�-�a�~*ԈAE�P6sI2�'�>m�e�O�UER�'��'"�꧊M�D�( { ��L��>~B8�%��y�D��3A��z��Ux�!�*>���T�Oz��Fx"�C5 :j)��ՐК5��1���B��Z�j��-3�%ZT�p��2T�U	�].([3Ī�H�^�|�D9Q�ѹ+���	���޵B��d��} 5Q?˓{
��S��;�A�s@���T�dY���5$�!���t\v)����z1� "�l�+o.]��4�v�|�T>��'����&�m���Ն�/YwhA9F+�18� ���'3��'�bb��m2�'kR+�(K���L�m��л�K�dI�p��#�hլ��D��8tA�C����OT�ʵ�LM�M�� �Ѥ4��jl� ���ݟ~/��S�i��1с���i�|#<����lZ�C��L!�g���6Q!/�u��z5�x��'��4�R7�A�b p�����*.��i�o!�G4q� �ǂ0<�@�8j6�DY�����4��Ē� N�uo�ݟ0�I����X��W灹�L���f\"3��O>���O|u��< ��,t�á4�P��Z���d�bb��P�j۾1kr(��m��HO�ܩ���*䔄v�Ҙ%J����G �|��ġ�+ݒx��M�ms@]K$�� |h�x���Ox�D�٦��	y�ԊO�tH���#E�ǢcFB����,�)�})��U�%2S�{[���ԁ
��p>	��i\&7M}�p���ٴ8Ʉl"��_� h��f�O|UxgæY�	؟�Ou^ ��'>�i�N!{�L^#&��y�+�	���� �>7����1q�ǐ�+�y;П��'��]cM�%��%�Z�ikc�I�{E��ش �d0b�m�(Wƽ��iE�� d⒗`δ���\c��{b��-b,�e�_�C�~���4p-B��IƟ�1*O�d�sӮ%Q�iAX����:��u���O���6���'��=�����Dr�fя@2\����$
���C�4������>
>=bL;��}�2Ḥ,k�$�'���'��x�� ��   c   Ĵ���	��Z�Jw)	  q��(3��H��R�
O�ظ2a$?����`��4ug��g"Y
d�+�܌�P_�*�yV�p�¤m��?	�'ΛFi���lL~��^�h���2�G�6*|m�!�C�s=�sI<���G�l�{H>�'��)p�鄺��ձ󬟦.j&Ry������۳�Y�Cl��ei�	���κ�-	&AGIvܬ�/I3_����@+LLp��@�rOZ�*c2�YJ>B��+e��)��>4W��ӂ��NB��U�-�׾'��k��|���8����'��d���<ƚ�����3ak��O������(O00�J>�S���l^PIɕʐ�a�r=#A���<1��*&B#<J� c^��3L �se6�ƍm���ɤ����^�,yB( �Ul���)��۷3}�F|�'�=�=�!�ސC�x��i��H���XH��-��I���,kD���4ܐ2BۇD\�	����t�b����I29��ɉ����2�ơeH����댱M��ʓd�h"<�/�	9Pj 0S��	J(h��j�q�m �ቜ_���C�'����Ħ��.a�H�!C����y��G�'�Z�'�<�we�^�����:
��+7���IG��2!Q��s�-�Z8"̺uD11�&XR#�O0��cB-�?)��/3���|�T���&5��]@���B�BT9(���a"��f�˓-xX�@ �P�,06�y�N$�9��@�O������H't��Ӏz�'kzmh�Ԙ''��Y���
 ��dzc,�,Y�i���#x!�٨# �  �"Of�'�ڌƀóv���!�E�i]�|H�C_�$��ŏ��ΨC��Q�b,i�A��W��f��q��%0�i&�OnТ'�W'�z%�"�����Pe��B$~#XE���_�Zb����ˡsI.�O��̱�G,,B��� <G>�A�}��N~Ԑ2"�S�Z��	� K�Z��6�&?kpEH���X�(=�d��iU�x�f7�'�~r���] ��W&�˅ub������*�O�x��Y�쳰C�j��ks�ƖP�X��'ֿ
;M�f@_?3�tTa���||hםN�'�H�Y�?�&�*�(л�@�{7���#��caQ��"VF�>��%�Ȇ~�,J�Bѭ)�8Lʕ���xy��y�#6)�F}BC�X���7g��%re4R0D`{�(�%b��A���'��u��'FH�R�xA�ءX���[ �~�A�74�d�S;��8��H̓R>��XvF�g
lc��	D�|��*WI��!��:�b܊^H�Z@�\.w�l9BbЫ)Ρ�e�o?���N�����7,ݶ.����GNN����������䓟:>�u�t�r��M���"j=�>=qG�-���1AĞ-�����(���{2g�&D#���5K0��P�M<\d� V޴�mq�D�:����5&�A�'[
 c�Z�w΢�)���0��o[[8�Qa�%v���aa�C�X����`d���:�����Q>��%�O��U��O�!d��=�Q&����1R�"�6DO���pE��GϘ�[��P�sI�$�- X�H@�&D^�|6If_��q˙�jێ�3&B�2��TA���ʰ��K�	��A-(h�ZP�̻D*ɋ�Q	n�����O?��<V"l��5CFC�E�%��L,�Kub�?]3n\q�A�&^���D�~�aቊv�|C��ӫ�ӂ��%����tZ�!��a_z�!�D�z5���g}�@*�7��N�h�p�;tڬ���^T���ɤ��ԴS��I��ܬ�-O'C[pb˼>s:�S���0qMP�9CKP0&���c�:gz��I�X��Hq�_�<�!�}P,�j�py�0eUF�vH��k�u�'����]�.H�~r���*$R(ԁ(8��B�O����2�RBD�RE�Sj��?!BR� +?��'~�D��ѻ+ĲL[ F�?+41k�'��Y)�E�B�S�����%�B�V��H�e	�($��҆nK��y�L� e8x��+o��x��ޜf��x)�e�  ��[b��6�hO����'�!7T�`��'�A��?yt���'D�ZD3$�Ü]E@� �8xC��D��R>��Z��\:�"�Q�E�Tb��z  Ke?����+��Rc5MT�`3s�>u�����P:���Dr�	a�Q7G>-�U�P�E4V��45I#�R�Z�rdS���� ���&��A`��)�,�孊=[tkbe2�Od[�%�:��Î��׀�iQ�/y���"����x���8=����"�Sm��PvM˲�hO �Ȏg��@��$X�;��4����=K3�+UB�8�y"e8'������7A(jU�R��ybB�
8%"�j�O���K¦��#���?zu�ңtS�4bе
*°�v��l�p����2�y�_D����#�b �ŏX���-a$)˰[8(Ј���O���WF���	B
f(��Ͽ���e�F��炑�r)b �ū Q�<b��R�])L��l��U��!�v�(qߕC��P� /?]���'P�Et�.�ɯ))��"�!]�|L~����=pN����-W���c�"זdf�B�>[y���'�<��Ap@+W�*p:��=yzR��S�? �I�V�_�� ��������?L���틾+>Q[t�V�N4�����T�Ӫ0�oET���+���wݘM�r0D�0J�O�1o�AA"���X�H% A��#v� `a3��!�T��e*Ԃ�>27�3mq��͒a�L���ޢT��pА#ـB�!�$Ύ&cНÁ �;q�~<ʗ��7z���P�Ɯ��c�G�z�"P��8�ԉ�!��8��'��ɡA�*�����5b��2�D�1;f��#~��X�@ d_�P*ƌZ�h��"���0FP�%�gƼ�a��&\O��Ƥ)5
�[#fN� |���b�	�YZ Z�M	Qm����7�8���!wܘ�a$�S3<u�H@�ɭ-�м��:D�����"s�� r�n�+K�����/ղ8� e�|���$	�l����RK��Of���\U�=Їe�Ύ�i�$�4A�!��Y99p:k��\�$��=Y%�"����G0T���a��[�TSy R�����$L���'���谯^;�h*4��<H�j���L�j�ʧ�Y�2����XX$����}�r�b���Uj�:
�4����'| ���8*jJ4�#�-.�%��}��K
nŲh�qd>#ᬠ9��<�������?y)�k )\��h
��.:dx0,&D� �G��t-�3B�
o�T�H ��!{�����W�>!���6�� �B(�'a�L�'h+�nۊLO�D	�i�I�QEY*m.!��*)7����K�.��1���F����>	�	�⪘3YF�t�P��� �,��',�I�VN�-mڄ����<&���xۓ����g$��R����l���`��Wn�MKH����f�;=©%&5Fr�{���.0���d��>b0�3�B;��'g�X����g��@�#��5`��ͷ�Ji�:�4as��#L��0�q�!@΄B� ��� b�GY9�S���L�& а�	&n���#_�b�e�T����~��w:X��FW���gj��qQ����'�^=@G,F ������� ��`K�+�B|�Zd 	�}E|�X����� ǬD�O}��D:2	�E�Eo�,�J1�b�i���XgfA�	�џ��'�@���ţw���i��3��Д~��`��߸
����h��!�E��d�|��t1�l_8�y�$%�������a��LY��3�HO�%p2��K��p��/^�C|�$�Q��?Y8�dO:����� m�B0�C:� l�N,�q�Z�PN��E�4kś9h�)-�3XL|�*Ο�9�G�'ڒ$�e�����D�ܴ^���30�À��4�`/nԬ�E�?�6h(O(�a3�3?���G��]�Љ��7���"����~­҇MK��ed�!MF|`D"	B�~��lç�l|15)jA���{��\�g�̝n����T���J��äK�(X�31Ҭyj�_������n�"��'���H��G�t
�kUU�@�F�B�+������.�'o�D\hԇ�Z���!�F[���P�<1��ۉ��`������h���;� H�0�Q�$m"Ё�`��6"=<O�ъ70H�\�C��I�� 36	��]+4P3ä�<���f�����eM��� �J�RFD�" -VT�!�ʗ����D�c�(pE��&��t��_D�F�+|O��P�&�$xMt �C�,��E*D�'D������f�U�6t�s�b͜3�fT:���7a\x��I���u¶��1�ʮZ�ȝ�>���-s% z���W^�P�wj�{s0!b*ſ,!�$�%	Ѭq�c�7����V�!���<򌂖��/9(�����!�*v�>���$�;ѹ��6L]!�D֗̸�©�0ڰX�FϦF!�$15���� L^�d��|x�䖒
�bG{���'�2�17o>Z������)��3�'�r�B�����8����q��% �'Va�N
$
�J����V�D�Y�J��p>M<y�g�{�@QDMP�rڊ�`���s�<��K�z�89�Ђ̏d����o�'0ў�'pL@)�a �-ov��c� ~54��ȓG��T+B�gT���D��]`@�x��)���`�$`�2��� A�f�hwG"D�蘧�.kX�]�/��a��)6���\����<]V�h4��I:�`�mU�r�H���=���b��h
�n
53��0!�Z�C!�$�]�0M�f_`"(1��HI�4!��\9zHE�%�!b�)�6'J>!�D:MFXXri͌vD(���S$ �!�� �h��D�JE�Zro�<S�Y	A"O\��CI&6��8�S#Ӟ=r-�"O������x%y���
bv��Ht"O�5YG���)�`�hkVт�"O�8)�FB�y����q��&?U���"O��F���HH�"M�%U@9��"O�ف��C1��uZ��ύ�ZLi�"O.u2�ר3��),�+(!��:完i�k�9 ��BL>q�!�d�b"��,��j��r�!��ݙF� ��Fl<.�h���<t�!򄚲r@pĊE�S�-���P�ǝ6fh!��#@ld���/�4ie�(b!����!�$��d�R a�?	Y(�#�}�!�d1z���)Թv4��!R�!���65�$Zg���t���]��!�Ѡu0�SgE1�)��Q&!��R�M�.����W e��@��$7d!�^�<�Ҥ[ԯ��j<B���X}e!򤒚�^�!�"K!/#�2D/H=O^!��XC<ѫ�[O���uI�dE!��F�b4���f�;:�}�dn��b9!�D�Q��}�ҬL?-t�
,X�T'!�=(E"8�`�],2��!�Ě.qB��G
4f����՚.�!��cl\�a���"��ɥ���<j!�ă/ 4��!:�(@	�
ߍ%<!�$����lǽ�0Hc�+({!��:7
j��tP0�ܐ�FL��3Z!�.ax��d�̍e�fm�f�[CJ!�RCarq;�G���.pAC�!�!򄇤:��$H�Mut	2Ta�4>!�����4�"d�9R�4mʣ[�]!!��H.p���s�مHԬ��e %f;!��>}�]����!\�(�� ��)!�$��]�ڜ� l��nŘ��&N�!��k��[��  ���!�q�!��.V P"��e �$��H$7�!�$To��A�D^��̹sk��B"O��
�L�_^� ���j�j؆"OL�R��>��e��e��1�6Xx�"O��S��l��04	_7z^���"O��2�*,Kͼ��G.T�zW�x��"OT��'�:#�`�/�"1�� �"O�}A��қyδ�R�)܈#"O��gE�O�< ��Ԫ(�S�"O�5$�� RМ!��A9���Ѣ"O`0�B8[�<� ������"O�cu���"ݺ���n(X�"O4yP�U��K��G�
�(�!ãR�R})uL@9#q`���*\j�Qf���
h�0K�'�4!�dԲ>���@O�cSN��cgB�32!�̖L,�I#1�r"����H&z!�X_�l�����T:P�P��B�!�����M��fH�	��?�!�$��N�6�5L�e�p�CD��z�!�/w�}�UK�+���0E	�~�!���?qV��rčQ)	�|��䑮Y�!�J�S�v��r��M~�� ^|�ݐ�'�Nh��H,NQ�A����ob�IR
�'��p�Ŋ��0�B��"�p�0
�'oީ�M߲L�L`�Ҷ	BZ�9�'��ݑ�`��J���R��\�O��R
�'���< Ш;@g�
E~d
��� 8E �n�2%P���ߪwm�%r"O$�á&�?A�2��H]F칊�"O�ȐQc��#
���@G��aEl�f"O��1��{�0��"F�i�����"O��yAO��Os!d$� }�z�y�"O0*4$��U�jT�A��b�h�"Oj�(t�SJd�U�f!K��|)�"Oܰ�n
�$p��ru��鰸�E"O�A÷\_R�Q B,>��G"O�E�sk�1n�(�棒�8.�%�"O��۶!/<l��$��&r��ՙ�"O�)�p!�AB�j�nLpx���'"O�H��E��.R0�!��2hyb�!t"OjdI#Q!c����DU;k�@є�xb���l��ك��'I`%(`�S�����+��u8С��`L�n�VC�	�Q�Ni�AD���l��1�_�(9xZ��[�D��cǖ�^;�D���|2E^�$��d(J�\�xq��6�Px��n���l t��Ѓ���/U�m�&oA�I�P Ó@�}��g9��곁��g�$��6��=h7�%�C'6O��Ѱoʦv���(�;�m"Fv�ꘪ���.f�BI�B	��HOH}
� �:�LTi�h)���Z�\� ���R���3�h��A9N���#5}bl�.!b�8C�VD��@�EBA;��R2 ׉7�z��,h�׋�d}ʁ(�T���o-��x�J����3�b>�#?q��R�!�L�+2�EcHex�-�;Ct8�&�Ԝb�xaR0�U�c��sćBo�'@�J�K��!Q29XQ�V)-��P1��D<���W |��5�-��c`k9
)83A'��X[����2�Rrb�^��bɂ$�C'R�Լ��J�6:P�a�vԽ��B�v�P�cS"�����������1"�\�d�R��D�:/�a��W!�z��^62�	�[8�q��S*E9�����ΓO�� ��S��кa��=7:�P�[���� ລ��Ov��@�$(J�ym ��	;�)��Ҧ��V噇M��]&��9�Ӂb����[�/�}�%��3�0*2�1!˼D�6R�$D}C@��E���*S��HɃ@T�)�%�bA�?i�0Q���|�D���>v,$����)ډnH�8;���>9�i�"�脀 ���	�j�R��&�6�P�2�7z��`�
�4Z@	A���O���ӑP�F%�4�T�oR���0�؞t<y���+���aF����7'#}h�CT�-�ġ���$���Ɣj�Aa$����'��D�� � ���*Z��m��tQ�&(��e�����^�%Q���D� �*��Z���{����Tj�Od-�Mz�������z_"�1�A���AC�-��-��袏>��M@�Z]�ܴȐ�'�YK���Bc@=V�(( uj�d��cȱm��!eퟠFH��#�	�\ٖܙ�L(\� |���_�v��e�'�B�`�咴+���D�;n�vH��a��&�V�Ke.�&d|t���a�/��)�������'td���ă
�t��+L�ux�҄��#�a{2΀+_�����J�G��pçS�Bh
��S//:|щ'�$��^u�6��>�� ����	/.x�`0�#�Ug�bP�)������Ql�4�6�(���$�V�[�Q):��] �f��1L�
�-[zb��ϕ.%�ܡh��Y!r��ܰ��Ot(K�|�8=.�O�=�B�Q>�)���-�dA�K�*��Y�닒8��ڶ@$Z2�<�F��ا�H5^��! @$ ��@:�[e~B"���{b덅F����d�ف@���M�6�x*�X�
ވ=�>9��"�X�S��Phų.�����O9���+��K����X��p򳈐�\]4�X]�lY�a�';�y��ԇ ��t���3:2�I5��6�j�s�B���-���X�*��Q�����'�(=�B?�raKK&?�n1�咽.����*�PH�D���3C����9�� �-��17��'l���Q�����xBG�/�8H ŎJ��􉮰�I!?�J�a��	hҀ����d�e�˯4���#�)7W0�6�Zd?Q�';q���Ur�'0̤���LR�����+H�9ȑ+�<I��2/ ��(WΟ ��ҝP�.�'C�bC�i{��#��)a�ɹ6({x8��1Ϟ|��@ޕ��'��PZ�]�OTN��B�U�.^
-
ş���啮(�L��������Б�������a�D"T�$���&��%3��#�$	<P�$1���
�B�D{B�Y�A>L������$� Q$�t��Oh��P��-��=�|�C���2�z~fR����*�8�"ÏQ"K�4���oVE����6�	'��0��1}��j �M,`�V��',�(t dBƾ+����'�` C�S��\G��0>��n�@3�߾g��x[��䉚u^�,m� tr�+�9|���'��6m�*�@����6���E'ܪ,��!�6�ɿ���y�o�0+��X��i�y`cB�P��^?o�D��F =�ؙ���jn���s�^�?�`��+�?�fF��?����|�	��&N��!D��/��$H �x�K���K�H�/r^à��	:���<$N��V�duЧ�O#I�\�e�b��<�?�e��
8���D/2:�Qv���&ޭ�'&� \%� ��KNЩѷd�;c��E�M"Ș���:=�V�� F*q���t�Q&MRQo�w�� �����`<4��]}��r��',�	r�R9u�(��?��!�{���z)��J;g$,���ͬz�8�J%���^젵qbH�"|I�ͨc�S˦�V��2F�T>�Pߴh#|��T�Ry�1���?G�2ʗl�@�)�O	s�S�ԏ�{��50��w�DL�&"{��E���/.�����DԔ�?��*]6Yu�:��$*%;$�D���n�O��~��9�\�<�|ݫM�,�w(	�,����Sc`�`bק-��	S<T9�卨 �ӲF�H��'N�p{'"�"ݖ4��HP*W�L�R�!�v���h��۷,!����Y���Pk�'ޯF�|��'r�I�������4�q��Fd��O� k �T9n���E^I4p���O/ޘr���N6�p��ł����'�����k_�yp��)D@�DJ�LY�A�?��O˻��)��`	����0�8P�G1	)�a��
�:���;wO8Q	�o�?L��CFT����'��� ��`�MK�G^���A�;����?9vaϪlA��	�S�8Mt���U�d	��^��k�c̿(Ȯ��o��N۞����Y2x��&�-g�6��<_��!�WM���8w�-j0��1�;WkP@*��4?)g
%6.֡�P��Xg��A�t��?�cm��rڼ��瀘"��j�-'D��YWbm)�bF�
'f(jȋ
c�ԭ)��_8o�4�rF�T>�R�,�7UF>��l�j��/H�>���x�%Rv�C�	�,0j�#f��O���M%k����B�-}�ɋ 
V��	����4D,���ᐡ��'0 �P��4m�8���H3>4ÓZL�h�©��>�*���L� LZ��B`���TT�n�P���\�%o>" �)�@��
ߓ{�$�coȎ�>��V�J����'�4|��Z���u���y��ۍ{���rAz����B�s��=5��ȓ/��<�!��/^�r����S$�4�vcڣ]��<3��H�S��H�o'H�k�w�|8q��1m��Is�	{�l��	�'��}:�M�؊ݳƤJ".�J|Y�����I��p���
1/���t
K�;V��H �+�nu�����9"�,O$Y#s��<<��#$�1!�$ Ɨ1`:j=agJV�"3N�:$�Q�V|���36&d4+6�4|O��a�I8O����Fj�g�<;��܃�ĢoNrx
r&r\0�%�韺}�&ݼ6r��a
���"OT�ȃ�-`���a)�)�ܠ�D��|�8p��.XqO�S.� �EGy��:b���/��X5D^�m`�hW̟X�6	�� �!	���&��Oǌ�uFRm��B��"I)��ňD�� �eŒ	Pƅ�1I7�I(��� |����H0�J$�1̃O���1A�6k	���4��+��)ѭ!�,y`Э�)��T��l�jTz`g؄'�勀�1%/̐�B�V�G��LZtjL��?Q�����S�'���"�)-�*I8q�L�^�R�����?�v���Sg��q$�y��2�i�!2���+Ҥ��d��7��mQ�gc<l��>�ʟ�D�T�m�I�1��k��:,u����I$\���bP�V+ܡ�V�w�P� ӓ:k�f��FY2Qa��� c��[f��!F|1k�-5x2Nۙ%�.-��hO~��$��Mt|(�"�'wI�����$Y=*�RCA�#S��Or0t�%���F����b�/�1ڕ��dQj�o�9X��9�'��'��Ua�#�����nk�c�@�^d�z�L��e��2.@R����O��A�e]�>����c����SЩ���(��A_�� ���
�rD�������䊤+r�3Ll��Q�Zջ�	W�B�L�I:��Q�!EP�p(@Ą�촤�	5[���T9���A=uh��:�-ӋE�b���*ϦW��Q�n_Lx���p*ΤS���.R�:�O�*&O΄��Ag�"DRԨ��x��\�;�4s����i��'>x6$CO:f|A2k.+g,e���'��}�"d�#;hj���
�
�XL�O�x�T9�������>]p��`��U��jJ�������Kg��"=x��O /����X/�xE��O8yc�, t0�:Qc���!���FM�DũZ��-:C�1��3����(D
�*ݧS3Vu0FJ�(��!�_�0��D*���O(I��%Z!l#؄S�E^�[��0$D��آ�2�=�O4�i'�,[Qи���QDv��9�I�6B@̰�>�w��fy���,b!�刺#�
�2_C �#��5@�&Lc�YF�<�IT�1�apVc�,�f�9'��ND�/O���a�U�@����LNjMp���.3/��'���Z��T�]jfC�.!��뉛%!���T�[(Dx@�GcJ�,:ρ+B���! 5;p&p�P�O\h���.A��؃7��|�?i�F )�NL˴��$ ��}Yq` z�:r��:4M�v� I��jK��$ Γ���L� pp�(Mi��hB$�|ӈ���"�p?1��;l� 8r��>e��8e-�3����B�Y8��׮���'Q(��W�OV���;+n�-3���)��$�!��b%��+t6Sǖ�&��ҁ��Hހ��y��	Lր�Bo�q�l�k6��]�H��`U�j�d�&[qXI��O9JuA�I$\O�����C���ye���� L�h"��E�itR9G3P�ZR�i�D�#��Q7a�@(�`��
������2tðU�1��!0���ϭ^��	�!��	��@�=�n�`rd	�!X*#=!D����6|a��لHXƝ�%L/T:�{%�'ڽ*�.ו��s�HX}��i��͋Rmr\�$�'��"��q�1�F�b�>!�ë�4��p{æ;�Oޱ��D�:e�����8g��0(���pt�k�'�1OƴC�Eͨg��8i@�QM4�q�S�;w)�7澸�C�K�]����R';�3"�sg�+~���1�>n���	""�,�$�B�j�	1�V�i���"N��0jʍtS$'?�d0��ZP!v�Ϛp�xy������$h�K�օ��Ë$W�2sp�s�X��ϵ`|s�jJ�|et�؃H��N�]����qԆA�D^�`�n��)Z�E�f�Ce$�����I�Z c&���`Y'71.�(!LʟdOI" Ҷ��?ٲIђ�6���Ȇ�U��L��8M����f�*8lIZ��$�p>YBK9�ưK@��0�����X�'���XG&�<҉$>��F�L0j_0]D��<
�LV�+D�ċFH�5]��L��!>p~�J�ͧ<A�I�p��;4#Lu~��	�����Y ��B��,$;!��Y35��!%��jR���$m�����O��CA� �P��qO���$߇~�6���L)HVx]��O��J�#M�9��1{Q(��bĉ�:%��sV����p?A�Lt1"A���1<T�;肗������Ib��N`�%��VI.��R!h�k�<��M��?�� ���JX�A�n�<��۲�B��fǌ�H�6����B�<6�ҳW�0�f�Q�� ��R|�<a'��:��5���\�
��<��Px�<f
P�7�S ��#��,�FL_N�<�EL��%=��YQn[,� ��u�<�cүb.0q*�]$B��OYt�<YT��Āh 猐5W"�z�)OV�<q�F��v�D�)�j�R�@sbXz�<	C��l��P���u���m^�<Y�X*BS�#� {�4���`�<�.� XR�Xj0��IZ��*E �\�<i���4��]sQ�O�P���V��[�<9�d�4u�<��-�}�ڔ�C	S�<��\L@∊Wǐ�O��=��L�<���U�9�@臞G{&���M}�<A ��[���!��EC��MU�<!���t�~t�D�ֻ	��XƯ�F�<�7BL-5n���&�! !��kA(�C�<A���JVdEb˒ kp$�GkC�<I��/oބ
��ނ,R4cV�A�<���� Qlq���cE�:�A�B�<���@��t�Sd��8���IC%x�<�����$��b�,Ȭw|(!��q�<�� [x{<�'�Q�(��#��m�<��N��O ��������"u��g�<ђ��l��xis�]�V@B�ɘl�<�c�i�Ys��
�Y��y�Gr�<�pˊ�8�|�`�˗�.��=Q���H�<���>�����oK�x�,�GVL�<�o�]��1��]�e&as�
F�<��)��fo��� #�B�^1��B�<��(
Z�Ar�?Q񺔨S��<��G�-/�$��c�7aH���y�<)���&��c�-D<A�c��q�<��kڗc�]sbD��c�|0`��	k�<��ߡPU,���d�te�e�<9Bh���  �D��5�p!s�F�<��Ĥ:�Xxd˂�-�9�P��F�<�+�<X2�-�����2�;"�[�<1	T�@�$��ĒT�n��%��V�<�%D��2�}�BC<(��qH�S�<� �� ^�]��a�%a�k#�\�e"O�e�� \4:,zcF� .1т"O��"��1tY$�ZY��aF�}�<)�Ʌ]�0�x+��|4v!6�Tv�<����[/ h��S�`�d��u�<�T��<�%���X��9Y�A q�<	����{z��*��u?���v�@x�<9�(�^[�ځC
u?�)
p�Uw�<��ŏA:xA{�nԭX%&�G�<�U��) 9!�I[�3���F�C�<sf�:k4�����8(��e��l~�<���C$Q��H!r��rP-[c�H}�<�`�;�����V�
P�f�_v�<IA��b�Lpy&��=^L4a�ufCr�<Ag�U�}�$tN��H7�t�q��V�<Ie�D/����iҋ�py��lR�<��;��5)cFl �H��K�<!�A�:
���/�=.�ᘶ�P�<��a[Iq��+bgζ)j�I�CQ�<IQj@�4�T-�ܴC��7gFJ�<�&T�;3�rì&��M
'��\�<9g&\�8���d��Fn�}	��p�<�ѠӮL�F,Qɒ�3ԬH�`d	p�<��@�$j�H�;|QX��Nf�<���r��1��6�0Mx���d�<Q�� 6���*��ŲI�l���F�<�֧�4�|���jJ$p���S��C�<�"�74�&@`4��;�pA�[�<aG,�a��|�&�ܷ}�����X�<�caҪ���iwiԞ5�"��l�<��^�X7V=� /cǘ�1��f�<a�ǂz920��-�.�ʑi@&~�<���jP~� �K��7����S�<	�M�-Ґ���G
%N4��
]y�<���ڎ)����c�I�nл�N�<�ԣ�Lq��{�Ä�~�{%�A�<1�`�3i ��.�{����Gc�Q<���s �yA����Իcd`���ȓk~J�Z��U�N��c�
\o~���	R�'���0mR$�L<���>�@ܑ	�'��<37A[�(g�H��F�A��p�'5�I�A��?z�,q��ID�d@!��'ڶhxQ��Ly�#M�+*���'ֈke!�"X��^��Y�'�lj���b�R} 4(��lh\�
�'P���) `
 TN��s`��
�'|pq�j�.F%�B��O��p�	�'4�k�#�K���b"O
[�d�'~R�pg�E�k��9�dK�@��4��'�r�q�޻0(���4���'4T��E-_ȾBc)uUZ���'��\�7�J�j%� ����d�d��'�&����"q75�� �&3\D�r�'qd�1*F3P�H���Ǐw~�!�'�AaS \2y( 0V*Ÿp�x�'�̑5��d^.�s5l�R|�C�'��,`e�A�V@:�4ł�X�f$:�'��d�d����|�t���'�.���Ϙ3��m��菱 O.��	�'\�,�"���{�f��bd�D	�'!m��dº�j��N��U���'��L��V0d˶pXCe�O�:��'��ёj�i�6�q2KÌI��� �'��-���MA��a儌?I@Nl���� ��aw-J1�h��K�)CuX1b�"O�`��/ޮ�Ї�)\�m�"Ob����%G�T�ɒ 0C����"O����	�!����0I8���"O�k�̟2��5��m�//(Uh1"OF�D�T�g��i��܆LZ�	E"O@×���` �M�|�$�"O�-�תE-I��ؠG�0[B�8��"O���t�	P�X�l�*E$|��"O��R���=\������C�c� R"O�Rr�B�҄�ٌ7�v�9�"O\YRv⌭:^|��V��=���A"O�H��^�����LHd�*�9r"O\eP���� �^�^��\��"OnT+��19�̤A+Y�t���)�"O��`�ܺD�H�*d
ݽ_�\�c�"O^|��	=Z�x��P���q���R�"O.PZ a�

8���DJI5VE���Q"Oh�Rπ]g��*	�,z��TAU"OF�:��J�Z�V
&�^�A"OhE2�(Wc@�$!���z���"Ov	h��::ʨ@@ F3K��2!"O���iD?J��4.ǩ ��+�"O|2�Dոr1�)eK��>��0�T"O�a�F�� ���w��4�X�z�"O�d:��)X�%k׫7;>N�[�"O�xQ�K՝Q�61�EM
�s$0�%"O֤3�)�7hBF`#���"ԛ�"O��H��()���0	��#0"O�l���H6,�i��·��%P�"O���Dُvf}!嘚u�N���"O�U2Gc��\��%�	 l�e�A"O�k�
Q'\��9Ra��"O\A���D�C��{� ��t<�q"O�q�BCXz������Z,�"O�	i���l��  ��W|}Y "O�ѫ���g���i�j�/,
��ґ"OZ�C�NM�fWH���F�&��Ȳ�"O�`�C�qڵ�"���\6A��"O��`!�8^�L�S��CH� �2�"O�Y�Jؠ]��� ���Q�@ ӧ"O&�C��S'ȹx5�>��D�!�W�/�J쀑ʏ� �l�y.(E�!�`J�8a���S���1L�v!�dJ.w@F8*����&/�E��,��/�!��V>��x��D�6!԰�$A� �!�D Bi�ݻ4�_؝�*��!��Y
�V���	�$���ՈN	d�!�d�)%�ؑ�B� A����!�]I>!�D�OF��cV �$"ζRq ��!�$8]!J��R���Y�	K"�!�dN<r�l����[;���Ys/\<C�!��.o*챔I������ �#!�Ҋ(uN(��GA�*��݂,��=Ǡ��T�.$�0�	$IX�����=Uv*d皹Qu�Aa��a�2�ȓS�\]:�&�S{N՚	^�W�|��M2�[���d�*�:��ߴp������]�JǛ6}&Ų�!2�6��ȓ���"�9��<��lM���|��+np�j�kA-N��5��oM�\S*4�ȓo��8(�*���DP`�I�"g$����`�Li�-�3)$�u`����u��ɇȓhX�!!�d�)T�P��Ĕ5Q9\��S�? Is2� A�|����[-��}Q�"OX�Bi��^�ȂÖ>��=��"OZ�b����Z���a��_�)J�"OX�є�K�� ��V���x�"O�p�@_� |�ړ+Ղ&-c�"O���dI<4-N�+�*ݍ\�*��"O���ď0N�Xj1*�`�^Q2�"OΑ�N����MHDGY�8۶U��"O�l�����;�8)Z���96��Y��"O:��C,��Я���\+�oYj�<���[�|��� ��6D 8��aTh�<�e������E� �~�ڡ�N�<���"pi�D�q��%:��8ڷ/�H�<�H8ar��p����!� g�`�<9��8F��k��$g�"	�À`�<��0z��0��!���E��w�<9a#r���
&T)h���t�<�Sꅵ�&;$f:w)8���s�<�� J�V1&$!� ^<��K�"�m�<� "w�4��K������Ll�<�[.ъEA���)�@X3T�i�<�խM>%�����)OҘ�C�h�<�u�Hx2F�QmK�G��a۰�e�<�S+�{�(���C�}��Q�Ôj�<�+�H� ٗ�N�w��(�G�a�<��ڃB=Ȕ"`�;WjD��][�<�3-�N� kq� %��%��^�<��m�>f��[#�@"dj�0b��@�<v�.=�&��W��3*D��g��R�<����*C-���P���lX�G�K�<I�
�F�J����֘�����BD�<q�#	�s18�&׿A���� ��~�<A� �6������Q8.�P�"�N|�<�Ul̾/�l�ѓh�2hH�P"'�]�<5�V���xx��2x���A�^�<�b�Q=iR ���M�+Hc�Xh�EU]�<i�`ƹfq��ɵ'��N���$�Z�<��k�596�����#r1�l�0��_�<I7Ș�%��Ө�N4�z�g�\�<�"lZ�<��ik��I�4arn�X�<Afޤ��;c#�pb^��[dC䉒�u���k���RC�+�B�Ɍg��4zgj��c6BL��n��%B�	"^"۶oC���%��h@�dO�C�I*Y�"(�b����St���P;�B�	 v#���Q)��XP.Þq�B�ɫ@�0P�Af��pAV�E�PX�B�II$Z1P��B�I�h��Ύs$�C��~�&严�Զ\b��J7k��C��^�H�KE��3������*G�fB�I�!=�i� �JH���2��@�-w�C�I�z�n(I�d�� KWC�%�xC�I %vp��[�o�D�ۓ��W�B�I�eh�����Ou6rɈ�� �rB�	�x�B�R�m?u	|X��K �V)ZB䉠��T�s�XM)X�a�Á�yR@B�ɠX�܉���0&q"�yr�߈FJ�B��P�&I�4��0g �{DN�4d�C�	���	#0�جH��aA&�_�QtC�I6u��X�D�	�rA��K��LC�I{p�A�$E��p�z�x�C�� 
�j ��MK�%E2E2D��
C����Ea�K;dʅ��'��^N�B䉕.)�R&+��j3�U=�B�)� *i�2��&?�6�Δr~�q"O��f*��&0� -�`�x��"OFA9�� �%�BК��(R�%��"OJ4�5k�9Nz����,Y��H:5"OdTX�j]3p���ȡc��x�$�R"O����B[�s��L���X��	`�"O
��@�;qr
�[�@9��X�f"O�a��Ť&춍)©��^���W"Oڌ8D���/���AӔ&�B�"OX�KW�%W|@YEoP�c�����"OXp�UN�8^X�pS�W^���"ONM@$dǶN9D��ƫ�7W���/�!�DUB�XB�
\�\�n��A_�6�!�$�4.���3�b�8�0�D�!z!�䎓Y��<�ǋD>�pi���?_!��'�r�PT��'1���8�- �x�!�$��4���o)��J��q��ճ/9!�[-zV�=b�gJ>�x4i�j��-!��RQ�u��� ,�PZ�
Vi!���*e�Ш#�H=S�"(�*�*]!��c� @Z�+�� �d��@D!�Mq����� ���s�9*!�V�LհU�e%V5�  H����!�Vz"H��ƹ+%n�(S�!�d��w�Փ4N�T| ��E��=|�!�^/C���`Ǵ����[�Ucl�[�'x�*�e @x\����E�p��'��)��LP/l˶�(r��6F�h	��'|�r�l&R�<�:1��>�A�'8^���"ezx8R��!6�zp��'N��(�lE�f��cA�X�����'�.m���� �I� ��^M��h
�'Ċ���c�9��=!A�ȆOZr	��'W��B���G
<�AP��O����'�d�)�$O�TUC��ךJ��m;�'34�A�c�-O���fJ�o� ��'�8���J���u���Q�z~1�'�BY �*��EB�\v��>r\ �@�'j�D۔ř�2�H�1�]�}[��]�H�c�$ψX)t�����ژ��%��tr� �95@<ɷ�_ 	n4��9ô����L�+���3�Fnܘ�D{��'�
�P��I0g.l:qL N��h
�'��8��p�ܬh·��а��']�Ta�.W6~���S$�Z>Fs�Ш�'>Ȱ��*
�i�J��-�05��|���a@��0jIp�Sv�O>�>T��	j��j=
a�gcM�?� �3��	Np���z<!j��O�Ԑ�v'2L@�`L}�<Y�Tr��)�c�+7q���}�<9s��zTvPYEkȤKվ�@5J�w�<Ad��.�b����F���a��u�'say��:_(ؙU��.B{�A��?�'y�0��A�"0�D�#j��/LtI�'�J��LYT���"HX�pw�5��'�ZH7>,��|�%�epA �'Dў"~��C�
i[�=���@�����j�<���].� ݒ��
:��r��<��ѻ?����Ν�t�Ĵq�C�y�<��g��[������P���ᡱDs�<��Oգ� ,�з@C�p�b�Jm�<�3"L�n�V����_�u����D�<w藏)-HF'#^0���*
�<�G��k��A��h +�a�w�<� �� ��6
4�

QS�"O Ȕ���=p�@R��9bP�"O�3� E	mʞ ���9薙�"O>"��;�,z��&#�B}:�"OUKF��3d�ܣ��q#|h�#"O&���[�{g��i�ću!
�J"O ��u!E�%8|2r�R&kbL�"O�	�����r�a�,Y��"On��a.R6#h���?G|���"O��3W&�"���"S�I�H�Hx�`"Ob�8F�P�D�nL�0i�l�vT("O ��B�~�$ ��I��4��'��ɞa$�a� ߇9	 ah4C� I}�B��<J|��ckX��0f�� X�B�I�\'\0'�E;>��H��!��L)<B�I2\���u�'3��1��P( �B�	�t����j�-D�nH�!e_��B�!�µ��O2s88�#�@v/dC�I>o��tsC!�)pV1�&R+=2C�	}��!����@�T�ۣ��Y�B�	����D
Ag�z�H D9�B��+R6�0����������:u�B��&8��0&f�mO�E�$&=4�BB�	�`<F�0u=73��i�fW'pS$B�	�l}4��L-v�X���|�,B�ɋdZ=Q�V55����E.F�r�<C䉜66�c ��LR�����îF��C��t�
p"�0P��5m��-��#<q���?��ƚ8I �DC�n�� Iam8D�����8`�� )��ϋ �����4D� �ƌ�;�F��t� b>���ť2D����ph��	N�<�H��Bc^��y�ôdA�AEH?	�X�傎�y�/�e��y9��Uj*��A�:�?��'�dH��S�2 ��;
N!�'O�|{���^�*�ag�7{v�'Q���!�
�X&�l��H<n�ܭ#�'0�C!! �>=٥f�e� ��'D
��c�-�9�C\�F�.�z�'i�)��*N�V�(r�ɼg��4
�'�0iP� ��
̎���I�83}Y�	�'��h��f�oJ�hA�J=#?Z� �'n���.�p�la�Q��,����'�d�r��l���1#��U��*�'W��(��0d�l(#!�ÀV$���'��)����:<��ga%VT(�;�'��X��
�!wr�i� ŏT��hR�'�&�����%f� Qඏ��_\.�`�'����t�6%q�%��ݸG�\�q�'���"�K/P]�S@N3�|E�'~tٓ�A 7r�B�C�/�)
�.`0�'}(���܊AP���,��Vb(:�'�RRa
E�_�]��&�x���
�'��
��	9Aʔ�����:���'F�T9��,t�8�(���0dLX�'0��*�M�6  ({��؈����
�'����Gj�4�|�5i��pT
�'jL�1�/��t�)�J��/���	�')���D�������K��2x�!K	�'�8A�Oxh�� 0'g(�
	�'��4���\����hVN[�'������@�5�3B@�Zq4��'G�S)] #�z�{c��:!̂e�'e�E��
$E�g�عE^( ���� �|�(�:F�U�Q�(k4�I"OJ@����xKT���n-Q�e��"O�MH%e�
e|Z��(L"e5�"O��f��'#���V��F8���"O(��R�!$@&3d,äMN�yR&"Op��D�O��ɨ��#�t�a"O�Ue��o{��K�k�`L�@�"Oʍ�$C
�U��(�i�"�NUYr"O���!��';^9��iL����"Od	Ѐ'����ѓƭ!���%"O�hq�oC.�"С4�G�B�na�"OBm�d
ʣ2��P%	�W���:u"O�)��ó"ԂIr���;��t�0"O�5���r��Px6����("�"O2���_���
V�V6��D"O�K#H�B�X5���7�܁
�"O�D9QV�q��\�-�2r12p"O�P�)ҬAm�,��끵M*��"ODpX���8x6X��G�"��"OT�J�EE�(��#[�\��E��"Ot�Z3@��M{ ��D�-!xUP"O�L���{�~�2po߮Ou��hQ"O���%�8 ����k�k�@�"O0�Ѳ�5.M��q�k�/
n����Is���)I�D�T���/�+����o	i�!���~�ze*g���r9S.	C�!��3���B� dKv1�@ԃ:�!�9.c����X<`H"!��K{!�D�'D6�hՎT� �tKѤ��k!�D����X��-�-��'� pC!�$W�b2��5��ZJ6qcJ��|:!�$Æ4�ȴ�/�<���΁~5!�$ 0<8��h�<BYU-��w@!�DĻxx4ۣ�I/~\����T=!�V���32�Mv�%�
q�!�D����:�J^�|r���)��V\!򄆆0W "0��4j�;Bu��'Q�zr����h�������4��'���e@�w�x�3iI�~�v�
�'�xAR%�+/�XJB U��2�)
�'v$,��G�J�� \�
:ڡ*�'�:�#��
"������l���ʓo�z x�� �����'3I��5�ȓTr�#�!��JY�Q&ӯ?kf��!u"�3�K?> ]S �-�l��=WT<P5/P2�R��1�^6�
U��m根I�&�V��t!�ڂ�dQ��Q��8�`�pD�a��;.�4!�ȓS �Y���:`� �XD��=�tч�!m<H�鑸?ud�)b	�NI���O�v԰TC@)�XxQ"K�*���g�j��DB�45 �B��S�Z����f����������s�b�7'.�ȓ8?��؇c�;x��Y��H2;h���W���ǉ�9I�h@ք��B�(x����!b2d��:1��^� ���y��,J�lq�pkӥ��$Ņȓb�Xy*��F� �
xx�Ŕ,Âфȓ>�8ay��ע}P(شF�
'Z8��x줻 㑽Y�x6)I�'����|KC�Q&r����7C|֙��.:0P�bH�h��4�pÛ1�ܨ�ȓ2chI	t�������:μ���r��Jqĉ�y!Lu5����8���S�? �,��*\+��!�m��"O �����������p�e��"O�Yi���xF� R�À3�B`;�"O� i�J�q@jX��E�̒�e"O�1Ie �r�� ��d ��I�g"O�51F�@0sQ������Sf�6#�!��ٳ:Ά9S�K2<��x�J5�!�":�	!���F[��q���!� 1s��`aFLEG:�:Uʂ�(�!�dTqѠ,���� ��A%��s�!������P쟍V�ة�TIZ�L�!�ă�p�z�P2ꟈu�|{vM��3M!��҂5$HfO�#xVe鵌ۺ,!� N2���G	�&t�u�U�!�\�v��I�惃*fd0Y֊�%k!�"*hIf��,m�l�"w�!򤇽F�}c!�"`e����G�!!�$%s�<��˽zE�(����P�!�D�ֺ}�H	�m�����
�!�D�	~0����'~u����E�A�!�"��<!��?HA���"=!�$�8_�թE�_�%<�`3�CK�Z!���*f�,�!BGQ�Y�9h^0P!��U���䛐k$T����?4!�C Fc������!Y�34	�8%!�dP�p)t�+���&}�dC��/=!�D$Pv�X!�+Y��X�B	˸CI!�͇�)�'�D��)8Q��[H!�L�	1�L�*[����"Gi�B:!��%#5:0%Ϝ/:܉)iҭs)!��):�p�RL�5q�PZV�(!�ϕG%"\�a�/cbҥ�A� �:�!�O���E����6&Fq��F�(#�!�Ę�xw�lZF��>���E�v!�$K~�hѡ�C�t�F�F�E[!�D�g�l�z�m�%_�xaܴb!�;O�Q%�>j��8@��Y�D�!�$E1V�{�	ܻx����v��&F�!��G'��)�j�
�(�vF 9�!��� c�&���a2[/\ i䮎w�!��M��p!Y���7,NM� �x�!�d�A2�����.T���M���!�D��������?i�ᩅ�٬3z!�B9>Q�k��$o,�9P�A$Yf!�d<m@����B)�pFNؘN!�D^5P��0cP��.=� ��֋YE!���ln��b��!rAjF��.�!��=Z{^����h�"q�ˊ\�!�d�G�
�"��@�E��`_�䫴"OMYbg��h��tG��?�5Z"O�=pSM�0�t�Y�&F�R8�q�"O�,�� Fp.1��>CZ�:&"O��Q�F�} 2�P�b�ޣ�]�!�$]�'Ϥ��`L��K�,&IU��!�$��,�|D�֋��(Dpip��O�k�!��X1bj��+�kN�eB�挲\�!�֋tL���Ȱ~ `�s#�7yu!��S��	��!a������3a!�ȓ{�f�e�,��\xB�S� !�������cGɚN�f�Pf�W!�DT`qda� ��
��!H�eI!��� 6]S������FY�O4!��4?!��+q"КC�����R�!���w^����b�y`P�]I�!�� $����|A Ij_�0��d"O@U� �ne"$`�nϙ�m['"O�p�ř�������*rʙC"O���G�$�`���LU�-����"O��3��le�: �@,�Qa�"O>tA��[���BM3��"O��{�C�.$F�t�f��]͜��A"O�h�&�F f�R�q䉒��ʕ��"O��bgH�^����#O1HT��"Oм#wFؼ% A�$�١I��s"O�L���T�̄�S��#� �"Ol}�j�#�ֱu��dj4Q�D"O�҂$ŷFL��fYAS$бu"O� ���7R�@�@��I,�#v"OlM���H����h��U?���"O<Hr&�ѳ�TZBMF�l#@��E"O(��H�JV^����X�dp���"OJ�{E� ��S�K<+ꀫ�"Op��M�<1��1"PuDl�w"O@�9��ϜLu<�1� �76k�4��"O�܃�U1F[�E#Gb� r�)p�"O�i��#k>d�㎂*��pY�"OH9 Q�O�6��d��d��=�p"O�l#BD�9�� ����d!$��"OhP�^(Q�! �oL�\���
b"O4�� 58 �w�T-;�Duq"O�sk�% 	*8F���Zz�yhu"O�x���Q>��آ��R�-	A"O�>>�{�iQ�t�VQ�SIO�H#!�$��<�F!��Q;��LqP�M>
B!��� >\d%e�'�p1��6(!�$U�?�@���UDFD�$.]�D!��<44ؒ��x1*(B�� �!�[MӰH��K�1%�T*��̕�!�䏡-�X�ŉ�T�� �F�=�!�[=Ro���3��~a|i�JĐR!���%�L��F��bI�=�7C	�fJ!�DW�
��b�V2�I��(2�!�E��PT�g��p�������{�!�$���2=����_��[�b�3�!�c����Ѧ#�F��e�+A�!�dD�����d đ}�hFX
�!򄞈r�|`s��5S�X��QK�;'p!�Ą!��AuJG�i�h�
���SQ!��?��$1F	K*Nx�1�琚vL!�dTF�2�ya�L�s��<	���kG!�$��9pH,9⪅-7�j��;U[!��X�2e�Ǟ.|��!��(N!�
�!����ɦ�Pj���Y6!�$�,8�� F|OD�уK��u�!�d�GmV�'�u8ै�j�Q�!����H<e�̾.R9%K��s!��Ǫ;B�<o�ҭp�Si:���'>TũFj�SlL�2@H�G�P��'�P�(7�Ku3��#�(J�شq�'����_�+c�L��K�.4C��s�'XJMCǡ�
Z���A�> ��'����̵+�R��5"۪T��'j���@3W�ȱ3j(X݉	�'_�` ��!&h ��M>�d��'Ү��u�ˮ.�$�G�͕\�♣�'����2��4^�$S�A��+((�	�'��H�g��_~����# �л	�'��x��B/k$�=���o��%
��� l�Ef��=α�&(G)Kv��3"Ot�V��h�嫓�^�Ek�1�"O��E�Q�y���0�dThrtٶ"O��+b��3{خ�b�!؂px^I
"O��`$��:���11T`0��"O�9�pl��oh�@  �o7��cs"O	(R��R��9%��$^칅"OT�"Q�"ύ�g��E�!Z��:D����ҩI^lH�"!k�0��@�+D�����9!c�#&��7��4BҮ*D�X�P�⠝zU��`1,�{��%D�lP��I����K��
��%g#D�0��Κ!:P�|���Y�A
�X �* D��CF 4#�2q�Ƃ�/�ܑ5+"D��[T�s��R&lޙ_0���a�!D�4�DB�*F�P�(fe�x��e[��,D��
`�(��dp�A��\Z�yc�)D����.�/�(���MF[~u��(D��bD�ůAN�M+�!�>jg��`�+2D�EjXO��9`a��9�1��.D�`۠�օ(�@P���#tDp%D.D��r#�0ZͶ�Y��GD���0D���΅"k�nɱp�Y�|{4	$D��aJȡ$>�]��!�xXp�'D���`cʂ7깢3�ס��}��/D��,l�-z�*#8��2�@�8T;:B�;�"��r��ӂ;`�́
w4B�I�Z��\ٷ˖7ES>T�Wl�	&�@B�	�jhz��'�0bG�L[�F<��C�	?A7��A3A��nΰ(��%?�C�<�@�*��ݔ,���"����C䉠9~�=���Z=�����]	~xhC�I�D a8�	ښ bjd�F�ȶH�RC�
_��GM[ZR���nǹ^6FC�I�O��WHz0U�I3-D,���'�T(jT�L4�*4��ϖU�c�'��@��U��]�ӏJ�E�Z�
�'+�X�퀙y�$�:s�Y8�����'�B�J OǦKPhsl��8r�m�'Ѯ�����P��%�3G��+'Dk
�'	�ːmʵv߄ȡϙ�Yh�� �'I���6eO�h0�5���Oh�19�'t���M�"$\�����ЏNi*0�'(��uj͈h��ͻ�C�i�Z�'c��P��1f$D% 6.��E��'��	[�	ʹ9��Q�U�� [|HH�'b��+�j\+g_�hhP� �"�H�
�'��i4N�w,0�2�n���K�Q�<���	�K��|��m��>�ʬ��E�N�<�j�L���y��X!B&��C��Wb�<!E'J�&�b!��BH.��KC"f�<a%-_�"�3҃��)�`d�wM z�<����c���R�˕:t^*��w�<�c�H�K�dࢀ�2=,V\%\i!�$[44*���*A�Uj�L{�ʜ�:�!�$D�N��3�; D(���ԄU!�d�4>��TG�$&ڥX�(Z�W@!�E�* ���'D[=1���yW-�I�!��W�=l�R6FL�J>�1f���!��{�q�N�C��0�N+:!�$�+B{0Q��f��")� �VB�!���I��[�c4�c��9U!��OJ�0��#M���J�/��
	��yd"O�˷���g�B�1�E��� ��"O� ݋��9�DY�"B�4ǎ��C"O�T[1�_�<=�c�a�-0tRg"O���%OL!q�b��� E�"k��Pa"O*d��&�$m�@<��/aUlYڤ"Ou8�W-���f��e;�}��"O�-Jf�R�la��-�F�95"O��� �ay���F :�hr�"O�(R�GܖX,�;� ��"4���T"OJ���掰_N��`Хb#�l�Q*O"���#*�N\�(U�4��
�'-�26��@�̴hBY�C�h��	�'���!��#d �!h����A���'���"ӣ(�A��	�5�j�@�'�.��&`��(i����;����'�f�8�ꉳ`�n���� -��z�'��L��J	0��0p�I%�6� �'�@9�"��Y6���G�.f%
�'n�a�L�|�|	��T�"�>H��'�ґ��L̙�b��Ū^�cX~Is�'3A;�\�s:�U)��I7	1\
�'0���-eЭ��`\�)�b�I�'eE�m���v� c螊$�Q�'�@`�6E�T�ABFW�D=ܸ0�'���h�M[���P�Ѕ�.L�9	�'7����?w��oB�Y���Z�'b��	���UW�h�U��
��
�'H���'0��D)U�E(��j�'�.��[H��@LI��� ��&�y�+�:G�Ps��(H*&�Ӗ T.�y�bFOjd�bF�����Q0�yR�	5�t�c��?������1�y���?��a'�ΌD��A5�&�y���j2�b���4|������yBa�`j�����_�'fz�R��#�yb��z����e�. �̓���y�27�l�"4nɢ׊���L��yk6���K�h�]��D����?�y�D.o�֥,H��0a�#�y�Cݎ+lB��fۥMֆ�0�R5�yR�	7*�\m��)�?F��ٰdƫ�yb%)}����C #Q*x�'���yB�S�G�,<)G는j��a2�U�y�1qJ���
+[$ r���y�@"Z�^��%^Onֱ�a옃�yB��!�^|��IB�B	�����@.�y�y�1S�@���H�k^9�y҈�]xA˱��!>E�!@����y�#Һlh�d��,S�!���R���3�yr���
*�2oG�	�����.Ќ�y"E�{d�ʡ��UNy�Q���yrIbZR��F��~n�%)i��y���!	]��
��g���d��y�m�N��\Q��_���i��P��y�前Ȭjc��;,>jg���y"F� C���AW�C) ô��Vm���yo
�C_�5��+ĩ������y��S�7�.��E/E ���Y�a�?�y��.A��))@Б��	��y��R=�}�f�U2(N"�pk���y�(P���Q����ԡ"���y�J3Y7�!���ֵ^ʊ� "�*�yh�c���R��ȅM���1��y���E:��S L:A��S`�y"Ep���IFN�@�>��ꅲ�y
� @KW��#0z�i�Aҝ���k2"O�cgC�MW��zTkH'`ޢ0xg"OؘBdiǈ
���`u�I�4�8�"O�k�g�.T� 	��)*���"O U`�J�t���k����"OF�U��#����T%Ls��=(#"O��xEC	3*��T�M'P�2()�"O�����y��I�#f͕]���"O��DoЪ{D�,#3EEo	��(�"Ob̃t��q �cNڂ[BŨ�"O�Ux$�Q��0�!V�G���0"O�� �ƦnhB(��l$��08v"O~a� `V�q��x�A�;Xr1��"OD�)p��G_�Pht�ǣG�tS�"O�M�V�C�MҶe[�KFL��"O��ȅD~�f����l,D���2�FW<<�E�C�r0�fL!D��X�T�����Ɓn��Vj D�x���O/b��T
Fa>V��]rf� D�L 7��)`�ܝ#@)\��qW�!D�p�7�C��e�[;�d���>D��(��Ĭ5];�N�9�,D��F;D�����8�`��4��5RTbq&D��3t��1(9@x(V�N�Y�N�8��%D�T붣K=�,t"5�WH6�
S�%D��A�D��X��@s�BER(�y� $D��ɖL sl����t9(4`#D�8���r�	j�B #=�;�O?D��8t��F��pjgIʈv��)K?D�,�$A#��U�4�	� �xHn7D�|�s���}p*I�d� ߈(;b�2D�\��{-��s���'�"�hrM+D�D	���V
)AF!ՌqI��	�"(D�4��H��B�^)k~<)��>�B�	
z�X�#ӏ��C$�ɢc��C�
]0�"b_>6�P�	�Nf�B�	�Da�aꡦ�	g� !�c�#O�6B�ɳD���S�^�@�0OǔJbC�ɯh|,<x镡b�z��Ǚ' �C�IzH�U �ET�5�:����Y�0��B��l	|�
��ѭqF֝*eە`n�B�7=���6AF�/�΅JQ����C�	�G�\@�f*	0B��uc�U}{\C�	*μx�D�� j��3��!#�6C䉎~��iÂ�24�:�v,� �C�	�\̀�UdF.4�y�dT*�B�I0��DA`[�~0��B�@��	@���X�C��3t��	@/�F[<�+�*D��� aLE������,�P�`�(D����IC�J#�� $�B�H��'D��7� Z��Iic/Ę*�jYjc3D������1Mdiӥ�3g�R���?D��
�&X+ʥ{� �}R��=D�b�)w`kG�V��
2.D�83�,^�JDV #E�:���0a!&D�L����Mf8iRR�C!C`b2E%D��ˣ��M��	c]{u�� $&D��J��d�X��1��+6X�
Q0D�l�+�-q����4`�Y���/D�(�7��
L���%"�r�Q�:D��`���Gpܹ�a]�<�6qI#�6D� ��oQ�s���bǇ�8B�2��o9D�`+g#̐!��u��CO�>:����3D��#�$��*AhvML������7D�� *!9��r�b5Ate' z���"Or8�7��G0��R2f[vR|B�"O<��V�ss��*�e��"�P-�p"O>��q(L<Wa0!1T�J�C�
VLA�<�ը�(�|�2b
�w�No�!�dD6@F]���,E�x�Ä�E�!�U�XJH�:��v+j�y#ڭ�!�D�dm�xB�4/r�T��#�!�dI"<��pq�.ߌB�)��A��!�DNwtdx��� #��=y��d!�[�J��R�	��vΠ�@I�3f�!�$ GJ`/��|_�Ez�G�t�!�P�-����3J�L��e�< �!�d�_��!	Q��<1�A��ƍ�zp!�96�΁"(J���Z�Y!��9/| Y5���eԵ0UD�Tb!�DY�&xL�[��?cs,�WCQ1�!�VN�|�a�1b��a�q�e�!��y�vh3&D<S�����ڦt!�DO�.��{�A!^�Ɋ�'Ga!�D�(�����)^Z$��K�R!��/-�d��͛�@S�Lj���U�!��*pH�P�<{�N��$�B0�!��7߶�US�>�R���,V -F!�$�2/l����)c�"��ыͩ,3!�6w\�؃��L��$�!k�3�!�D��/�z!šƌY�`�C�;�!�D"P
DXW�BmѾ��5�ފ7�!�$�%&BH�����Y�2�;�.�w!�d�78"���GO�l9�'o"C!��-�lyr�E)��(�����!�d��|�V�Ұ�S=̌ÁɩaW!��PJ�m"RF��)\����
B!�d�!R(�{��_��}�!��9r"!��(!�,�� .�f����#�=8�!�d�6�n4��
�ΘQ5lG	3j!�	�Ёc# �a��e���T�!�d����tO�*-~��W��� �!�D�?j�D(	�뉜ªT�VO� �!��mۆ�hԂ\�%H�P�$$� m�!���!����׈^H�z�bdJ/th!���1L�p�B!.T}V&P ��ϟ|8!�䎕d��yQƈ�D^i�w`*
!�dM�'%�!�NY�);����.@/Q�!�H��`A���3h��ch�,�!�d�b:t�b��:���f�(U�!��e��	��1<B��̃w�!�d�?�����O�b�Yp��
;�!�$�(Y��@���"�n0�O/#!�PS�*Z���6��x�D�8gf!�d�VtJ$KBO�7���9�
�I!����U��ڢu�TT�@+��7t�8��J. D����U^�!�wǉ�1Lؘ�ȓLJ�	��D�;	�Ґ����Ԇȓ[]&���onT�H��d�u��J0A衮=~�t�g���@@�ȓ1�tX���_��]��c�Z��)��T =ze�) ]0la$�.�n��ȓ�I3�eM�ohJ���_��p��c���SJ�D��p�Ũ
�R��8qb���[�d���Nv��T�ȓl8lȪ"^bФcPK��p|���ȓZ"İ�̝�$�$���ғSN$�ȓl�a tF�)�>9��D��|���S�? 
"�dˁ[ؐ�Pn��W�0��"O�Ub���Xs�)q�?B��"O�
��:FB�𮄦P�I2�"O0�����jB&҂.��+߼%{a"O`�*T�Jx0 	��?S$�5Xs"O��K�0Qj��E��M��@�"O��2��"]��R�n�> �>�%"Or�9c7:e�msG��&o��y"O�!����!XXj&Кp٣�"O�D#4��.E����f]�4�2�;E"O�t{A/хo�T���^y����"O�ԩ^y/f0ӑ�W�!�"7��b�<AP��A$d�A� �Ws�YQL�t�<)�ƃ
]�PL8 G�x����[q�<�C�rR��gΈ`4�u)��k�<�fO�D>���t���;�]� jUB�<���@�	EJP��49�@E��� �<��c�0F�&y�ej�1[A�Y�B��`�<�ϕ2:���h�/		/J���B�<qN��s��}��m� ��D͂d�<i��X� �:��E~S(-�$"�;�y���yh�ਐ ѹaɒ���y�*Z�7��u�_�%~<�*�']��y2d�����0�ěN���K��y��I5n-1��8��R�O��y�"Q&��tP�d]�8:��g �y2G�l���@(�+q��X��I4�yR�Z�X�!���p�&���y�bRf8� 1��ŝ|Z�5탁�y"�)��mb��X�Q��rT�[��y�8+.��L� 욒a��y���#I�:�H�q|&� �����y�		6E�HA3'��z|�e���y�jV�XR��c��s͞p8"�_?�y�*�_���P_(�XVA�*�P|�'�(�iю��<@"愈�
�n���'9��p�Q�V��U�ą�VY2,��'T~����~$������Ѥ��'����T�
p�p �ƽيp�	�'f�	��'�8b�
d �%A�� ��':v���Aҳ>6�X����xQ�'����͂~���e3f9��"O�X�3fR�vּI�UJŀev�j "O�!��&:J�=���4"O��V��E����v:F��=2�"O��c��<W�V�5��s�H��"O4=��(U�0�)����Lt�$"O�q�dŗ�1�\)�pȚy�"ON���l�l�Nz��ڿz���"O~ �1��53�&-��L$<�A"O��P*��r��î���;r"O`�XB�]�?]���&�ٝ<�ЫC*O�@9��O�P�� �%%��x���'֥����0yx��
O�|J$��'�y�o$�I��b��)���'Oځ���V�����"�(Ե��'O|Q����?B�h�p*5I���s�'�`	��I�6PT�jU��sV�l�'d��FC/7��\XTB��q�h��'݀0�G�GjV�a��f�l���'��i��T�~�)���ؔzP���'�ra��ȧt ��G�Y5�	�'^Z�bmO��E�C gz!��'aT����%���	P=
������� ����b��*�>��'`�+g�04z�"O����$'R�(X"i'4�TDS�"O(XIфW,Y�����.�d"O�d*��0)Tur����#vt�"O�0P[��
���ޜ	k�IK"O�xrcc��P�r��g^v`��Y"O����ϡA� LX���%E^�dB%"O��8b(�M��D�G]��zA"O��^�N�*�Y�!B){�T��"OZ\$�!9&��;C���b�""O�u�ׅ. �6mS�����6�[�"O�4��gQ�����@K�1,�8���"O�؋0Hϭ`�.�������Q"�"O���#��&	��#���%�b�5"O����@��j�l��G2/��	9�"O�|В��9�؋�	Ɩ3��0�6"O<Xr��ٙ0�ZMX�.�d��!�"O>!p�F-'�\â�fh�E
v"O~9��nE Ē�{'��1�BpU"O�u�̙(�8��d�1;����u"O.msw�޺VY�H���T>pv�I�"OT9���=3�(�4c_	1_d��"O���c�'Z��EARj�#�"O��BA�C)n��4��=h�V��"O4��j���,�&*�!?�MY�"Oj��d�D�#����H��4#̍�p"O�s�K�?��%��.����"O.�sԅ�.F.���煈1֭@�"O&����ݏUD���g
�=��p%"O �P`��"f�Y !���-�Hh��"O�8��#n_�pC�B�;�� "Ot����Z4Z�(���� Hԁ"O&|��ӸN��]�4͚.=B�h�"O�(�2�J�0���U'.�*�"O�u�PjE�'��!v&�+[�T��"OjA�!J!8��u#�j^��QF"O�a���j\��� 
N��j�"OjMb���)\Rک�3���@?��c"O Ԙ�NE+e����"//:���"O�í
��Z�����~p����"O��B��]�R�t��z�ݪ�"Ox����
h���.˱JR�ѩ�"On��s`*c}�� "�G�Y>�t��"O���
_���H���970���"O�-��!�&s�v\�$�S���#�"OtpjA�V3��A�-ȏXh�k�"OZ��q���XD*���\]�blg�<��c\Sn]��fٿKp�ᑨ�d�<�6���B{�0@�`�9P'�-�t��a�<A�쑏@?���X�*�ƭ�CD�b�<9ǋ�j�&�����2!v
�����[�<�q�=�pR�¦g#di���V�<��c�1DUЍa�aC�6�ã*�x�<	U�ۊ�N��jV.N󪜫㆘I�<�@��Jm"a0��ʪj�&L���D�<�� �'f����N�t����Kx�<��4Y�����h߭.O��G#�w�<�K�H�v�1b����% 4@�Y�<Y׈өdj�m"b��3�(0Y��OS�<�Z�������|�ȷ�YL�<��.��UcJD��!<L	D��҈�F�<�Q]��H�����)���p�Bm�<d��V��R���?�:��լ�N�<��+�Q�Y��ʙ%XPf�H�<� ��fٽD�Fq*Q9�Ͱ�"O���F#�s����(Ò8TTC"OR�_>X�1�L�i���2�"O��
�-J�%�
�`#*"<s8�@�"O{�p�H�8� ��3Ȉ�����ȓ�D!����nh
=��Z�DІȓ;74�QB♬Z@,�E䔉�lA�ȓ;1j�R��C��2���XC����|�����>�R=��\�Q���ȓLiZ�;�N�1%��; �ٹ~�����7�,�+��I�*1j �7 L����t��m�O	#z�����4R��C剐%����dU�t����1��C䉊j�Lp��h"l�
�FCd��C�.BC:���e�Xp�悋p��C��7^���e�>�e	�aD4;�C�I���S�i��m�8�����JU�C�Ip�9�"ו7�"4+��_9�C�	��,��ba��	XNl�w��#2ʀC�ɮ���K&�@�=�@�:R�OXC�[$d4)�kG6��㨈�9��C�	u� A];!&<3��Э2$�B�I� ��Q�D�$�(�ր�3$��C�IVN�PA�1m^ <�5���a%fB�x-D���	*yR���Ě�Z�4B�	/��yR/��k��q�1d�rB�ɧ��e�QB3V�f�Q��\,~d�B�	�Z�*�YE ��9,��CY�OϴB䉎��Q���$S�@r�9t0�B�I|�t0R(S� ���5��C�	{}�x�ebM�D'�D����C�ɓ%��C`��K�6����S"O�	r2�\�I��\�U�W(\���"O
x*A�O�U��%�0�E7=��t�&"OΔ��_/!�4KE&x�9�"O2d�׬A?��Q��
�v�<�"ORK�LI����Z�NKW��)�w"OF�JB �7╺�oU'n�X�8�"OJ�)%�5wS�yi�B2f���S"O�Dŏ����ڑ�S�|Ǝ��"O�LX�Ne�l�#�A�?
�2�"OF�!.�jN�\���f"O��(7�b�~�B�J6aT��"OF(�ĂËh����@�ʸ"\�4X&"O\dJ�LУs
��5i�uFT�:"O�q��3L�*P˄�<@�f"OD�.��t�F|�ȡl��I��"OL�;Ǉ�)��M9�5��p�w"O���w�֣=�8�k��@�z� �P�"O��zׅm�u�ӧG�0�:��#"O<��q�1ʤ���Ab���G"O�P��V G��+E�sD�<��"ON1* ���h|��rW �T�@)�"O|�rL3U.(Zr$�=e��8p"O��2q���)g��R�(�%{�s"Ov�2i�&g��*sꎮP�A�'"O|5�Q��rv8*��EK��q�"O���6�]�)�>�X�AfT�|0�"O�ӵ�J�)�4IS��.GGj-��"OHj�b��1Sfp��/�/Mڧ"O�9���u�Ġ �*
>(�9�"Oа�(�� X���M�@�e"O2�0J�:o�v�ӡ&��G9h|w"O�����:%���j0��u��	�!"O� ~aC�YjJ�[��O�}ߐ)C"O��H!#Ҭk�Nao�1}O�-+��>D�4A�E�5�\� �H�cw���)>D��Sv�M�8ȩ�0��31,���*7D�Ӓ��J0��:6G����-4D��!J���8�q^N�l�a�g/D�P�`l��c`�hb��3PŠ	�eA!D���1��Ȗ�� B�<zپ��4D��
2F"1�4y҃�Â7ְa�D$D���3H�,�tx���U�P��U($D��:u��R�ꀐ���]+��9��$D��@��/���S�V�Z���e�<D�ࡡƀ��� ��Tv��I!.D���GO-Ngx�&��X�l�b�1D�,�a��E���L�P������*D����)݀�
<�UҺu̴] ӡ*D�<bFI�?~>t9��Q�;����*D�d"ф[*`��[�J8{tri��;D����ĝ�e��a0�ʜr9��6D��:Շ��o�:�) �ıtz���H/D��(���H��8���ޕ7b��iw�,D���� Z��4Sw�sh}K�)?D�t�S� `vr�R���H�1�$�"D��I�,/oY��x�O	�_-Ƥ���!D��	G�V�lz�U`bm�9%�� ��	:D��k�'��%����g�\��˂9D�xT��
���ģ^�č���6D�t(�Bы!�$�7�E�;˔-��3D��8a���P��N��(_P�p�,D�$H��H��d�+0&if<Kr�(D��ٱ=#�� G��p��s� !D�,��ߚ,�@�S�`��t��|0�� D�̫C%M�n���pC�V�Aٲ��*4D��XrL;��Y��@��~�p��0D�PQ	Ѫj�źBa�	.����@.D� C�PY�0"6Ǐ@S�9�4	9D�0 ��,]��Q#-J�9��4D��"���0�u{��@7L�	�J=D�q�
p`u��/j����FM<D���kB/B �ᢀZ�6@�%�;D��"�V<�4�&��_SV��ŉ:D�p�;��P���&k�Fa���=D�xЄ ۻ}N*,Ф!�67E2g7D��;��G�@94�g�M=��s�'D�d��M�VHbwi�3_����3*"D� Y6��H��3A��_� �2�G?D�|A��F>�P�&�8p����fA>D�h�6K�r�����$� 	9�D/D�����%=��!��Y�R*P�g!8D��҂��6�>]�pGԁi(qU�9D������h�v���h�?Q˰�R�<D�`���N�t��W��#Q@�05D���enL��7dT�HGĉ�3D�XG�ʡX� `�,MVQN��!'D�$�AJ���2���>��� D���A���##>��ID���-!
�C��u�j���ժcT(,ЭR3�C�I-�M4)��JtȰtA��n�C�ɯ1�bL�r,A�a���_�/�C�I�*P��V��;�e��'�A�C�	�.)d�1��
(�QSǣT�-nC��"(�,ܱ!䂋KﰡR�$R
P�C��,&�^ё�OQ�j�Q�tgP=z C�ɨ��$@u�N*/L�5��$
�C�)� �H2v��4.������ı_Y� �w"O�%fa-�.�i�*W�!S�T�"O�qHs���_�f��g�X9,��)�S"Of �a����bM\�6Üi@b"Op��s�-$��Q��k�/p�V�#"O8�ReGƴ9�8�6I*��ec$"O��P`���:r��#N��S�����"O�IԬ�4 �[`ҽKm`Đu"Oʉ)��,O@��ɶ�
=8�D0&"O�p��7V�B�H�V3e4��r"Op�I�/R�#"�;��M�	,�,�""Of�Q�hK.I���0�ꀕB*hؒ�"OT�å�/g|�K¯�,%`�b"O�ܢg"փ@��`3O
3^	�\��"O�i�E�0Q�-�nI>,	���@"O$����@�c���Q#ȃ3M����"OzT1�� 2\��R`M�(w7�L��"O�ir�GSy��= �l���p�"O�(8�-�hYZ%�H-$�3�"O��C�ǜ�<,��P��I�"0�YP�"O6ѸХ�,CP���dL̡�<)�"O�I�pa�h�	�@���&"O���/P�r��H
2 ��E�Q�"O��D�8��*��?_��	�"O6�
w" jq�0�o��S�PQ��"O���C��-Oƈ��C�>��b"O����Dd艦��	�)*�"Oh�Kb�"��a��+��oT|�A�"Oİ2K1%j�5�E�^�R8�"O@y��n�{9��I�,�2�ڣ"Oj����r7p��� � "O]xRF�!"�T �&�;~�)5"O� ˶�N�>�<���gh@(�S"OH���� ��&	s���	Uf�a"Oj�Z4kP�A�,u ��� 6*�$"O<j�QAnq@�gL��`S��2D�����z}K��.�J@��5D�T�AƑ�58��G��,��3� D��J��&X�zp�5�:�<��>D��bmnNʼ �O�t���R)D�$a��u��dk����ִ���N�<��CYu~W��E��1(��E�<i*=A�F t�����A�<� ˯-s��1,�"�|�1����<�7�R(�
4�B��&�"����Oy�<i���"S	�m���{�}Y�q�<��'óN�H @$P�T���q�<�5����uS�.��7=4 ��Tk�<�䨓	Ȩ��$iǪg�8�`"d�<a�@�>��n�A��6���y"
��`P����dQ&M����@��yrf�8L-�=�rH۝.I^p���?�y�d\���gC�)A�`k!�8�y2�_� LRYz��°.N��y+Y3: ��e���F}������y"�_�3	��2F��+%Ibl�'�y"�/%���AH�oJ����H��yHC�_�"��l��y&������y���I.�@��!U-���1���y�J<[��L0�O�"���Q`���y�	���x0З��6Y�-��y��)�t�2-�|Ҕ�����y��B��{i��m����p��.�y��U��#q��-\�`c���y
� Pp�ϋ�T�vZ�m��2M�h:�"O���2��
s���FQ�fC�1"O���dm��xW�P�bEeԒU30"O:xb�W�$�B١EH��0�"O�d����L	�ř���i�Yx`"O�5{��7 V��BE�1L�Ո�"OJ���Ɔ�ph�=�'�E?@<yh�"O��� Ӄs�$yU�ˋ3Dဵ"O��6�_�}VF� �ʏ.v ��Y�"O�L
�T�TU �IU�Z@���&"O�8�����Ď�r�	�s��l��"O�{O��K�f����ƙr!.���"O�]s�o�:'�{'(�_�qӶ"O�P�4�P=V�0�JgԈC]�=s1"OX���L�M?v���囤;J�p�U"O�9iSk��y{��0e�n28(�"O�:�i��5���ʧC�g�4��&"OҀ� * k�͞~�` 2"Ot��L�����@�
!2к��"O��;��� V��k���@��T��"Ov��5A�(]�HU�5G!��{V"O`��KZ]2�}SA�[�q��x�"OY7j�)@�zl�.h��3`"Oj�x�L"*��P*�4�xEe"O�}B��	2ʈ�`$�2^�x��P"O`t���J����k0��`��"O�BQǨ6��b4��X&�A{E"O���Ҁ3`��#�7]���"OTh(�#A+c!���B펁&�TL� "O��0�
Bu�iq!" x�F��G"O2%r��>\�.D�t�NQ�ڌ�f"O>A�DW�~8���g��.��]�"O�������*��D�M9�:pv"O�����#$��C�ۚ�&��U"Ox�q��Na\���ʻT@���"OJlxFۊfT9�^��`�P�"O���ūñ~�Y�3�%QWu�&"O�if�y� ����\�=;��"O���J��,{��B�vYj�8s"O��"6��8tc�mx�!ʨy���r"O���D� 5}5l|S1�T;-��)
$"O �VMՐCi�����&t�M1�"O6�A�S�r���c�Z0AZl�)�"O��[fk��鞄ۀ�>dLʼ�B"O�$	3MŚs�ZI�d���0�pʁ"O�(6��(?Qj��TF �%8uK�"OFy��� U�s�T�e{�"O`�6��#A@���C�ݻ~�
x(s"O�xRr��v����E<2J�h�W"O���脸 �̌ ��?#Eܨ�D"O� hd�=Jǐ����,>hpHe"OxD�.�+2I6Ma�Γk*���"O�ȩ�DW�F�P��B j�ɀ"OF����e��u2qX$� @"O��
��k�b��ԫd� ��"OXz�J��&#��`o
�)�F%�"O0<
�Q�F�H`�W�U���"O|@�0&0�^�aC��N��ó"O�Us ��{r>TR&(Y`�@"O�#����n�"B�<~T�a7"OL�Z�MV�m�vB"��I��л�"O��ؑ�r  �Sk��i86���"O�	2��_#~�P�a���  ��"On�#Q&��fּH�Щ�u�x�"O� 0�
4N�Dՙ7��C_�8�"O�q�ɍ/V��u�Ō\"dJ�"O`-y�@��(��px�j�%UMX {"O�U���3Y{N\��jƻ5�@l!�"O�A(#�ߋU�l!�E�{�l`"O4�Eߒ�����dc��!�"O�	T铋��T��$GJ uC�"Oj �I�(��q�p��9m,�D�"O�u+d��9-K�1ː�L&\C���"OB9j�Ǉ2;������BUa���"O�����{%h%��ү9>���"O
lx�#��-A"�HfК1>���1"O�y{�EO
b���"S2،i1S"O�xZB�.9�t)I��Ɗ~�-x�"Otarp�LC�ٻ'���?�D��"O�����ud� ��H���fę�"O�S�@�p�ur��_�`G�d)�"Oj��� 	������+1И��"O����5���Y�iBӠ"O�h��^@��f��AX�3�"Oܨ�KQ�v+�)�%���L��	 �"O�i*�R
' Az��ׅ��AC"O4�@�QD��I7'P1Ur��"O+�V)�B���T��ًpKGc�<	��[�ߦ����G4���DAG�<q"&��!�Q+�6	�Xc֩OD�<�#�Nh��d��x�X��V�<9$�ũx�:H
f���	UԄ8s�]�<1!N�8�� �pBU���d�P
�k�<1�Þ�!���a!!�s�9HG\�<����7�p��H�[�L9�hDX�<C�D֜�띄e4��B�V�<	)J�{�L�
��ԛ>��0uƄ~�<��㌂8, �.�>P������y�<I����i��m1�烄R���cDJN�<��G�F��=��bͷ)���8��B�<��N
�k5r�Qj�*)����@�x�<���ޛ$o4�h�آ2u,�x7h�u�<A`J '/�V���Y p��s�<y�$3�ބX�!<A�.Y���v�<����!G���#"�A>�%���o�<�dHٛ,@ԹAE�$? �s��S�<���15��p��]h�^���j�<�söF�| �6CV�A;�p�A}�<	�bH2<�ܒ�Ɛ!P@�I���b�<�k�O���@o�2/+&Ts6Oa�If8�0(���'`2E����4F�*�R;D��A��U�1[�͛��
PJ�
9D����#\�RM�ɃBת6�lZP*)��hO�Ӎ`niA꜒�l̀1�ڧ�nB�%�A����O0di:�[���%=wў���HO�,9���R �պc$Q�ƚ��!�$�0�n�XL
Fx�<Z@`^� �!�D�g�`Ч�<`�\��ѝo��{b�ڌJC���A�Q�@�y���!򤏾y���
D� �JGj�OjOH�I}�O֜��r��' � jh"O,	QgDL{q@��m�V벍�����?����O��� 7S����O5�̸�"O0a	�@H��V��0J~Θ`�6�d��(O�'��<2%b��g��L2D�/q�(]���� kF�f5�Y0��q��Fz��'��`��K�>$�� .A�4�t���'�Н��AI�g ���$ņ"cj�c�'�
� ��CG&���F�ِ�J� ��jd�'�qOd����J��|6���&�3T"O��q�	I7 �	d�� r�U��'�;���9*�r���0P������)=�$B�2u���Ж�ۖD�Ii
�Y
���5}��'��x�O�r������'&���ち6��a%Ï�ݶ��'�ʁ��	y}�ڡo����'��'�7�0§���C�{�	�J@r:h��$�#341O��{��?y���7Qve�L��UIfӎ8���A�F]��l,�T�P-v�<0
��
4� ��*�a$�فe����DC�q$���k$9��$ɆH� ؑ0�O*P' ��vls�'$�"}��G��y�'�F=R���p��Ա��B�I%tNсWh�.J�aZ!�W#w�VB��7|�9a2	��h̬�� bUL|����S�<1�g̑f��=pC䕯��zC�F�Ĵ��鉹�6����7J:�3G��}��I��HO�m�-�3��&Dç?� b���x�<ib�_<
T��;D��Y6����_m}�Mo�R6\�i>c�ޡU�dH�U��3���HS�!$�L���D�D`b�
��h�ƃ�K�<I��ӝ!B2};Tb[Pv�H�V+M�'�?!0��&��Y�Bk�G�`��!k?��l��0�S��P3<�y3I@tO!�B�I�q��'��fO�1�W�ɦ^�lB�	�52���͞"����� C�ɽ���]2u?�]�U��3��C��'�|+�X	T�*�K0�D�=~�C�'![��H�$r�y���B=�C�I	�fH! l6q��[㌎1n��C�	1kU$�4�bd�UA�4O��C�IL�8�쀩����6��bVB��П�z�@[';�N�˃�T�myb=���$D��5�4FMJD��'�Y���@G�!D�ȑ0I����xUC~�2��/?D��x�/#x6 ���F(
	�7.�>�޴]L�O�>yB�O�U�<�G��?N��k*D�X�W�E5%l8Y��G�*Qzvy�d�&�O��	>a����L�pۆ	�偕:<��B�	צ��fN:g�tX�&��$�Bt�Y}��'�F�(@�H'4o�{=��r"OL�"d �	�������A8%���i�L��	�	J6|�n� W�0TQ��R�U����6n��6��x�k}BiX"R�yr���z0��A#�y"�^0��-��C~l���b$��X�hʓ~��)�'4"U�b>��Q�]�b��XC��>W�r�X�5\O7�#��*l(Lsu
�(u���'D$m(X�@��	%A�����kI�f-��s��@1Z�c�h�O66�/ҧE���W?& ���K�,�xi͓��?y��	{��("D!g0D�����zy�HH`��H����H�˳��"����d��s}�'����*8HxQ�)Kt#P�2C�)��<��M;9�i��"C�`Mke�X�<�g�P�P��09�]��@Z�K�F݄�2��`'�+��1p�né:!DB�FZE��"�$7�=@w*��d0�ɞ��ID~J~�'�6e:�
�1}R�Գ�h�&s1v5ش�hO?7� �p���)$���������,dG�	}~��'N~�:�'�	�(-���Ź4̌�J
�'���ӖG�8<q�����-�M�
�'����b�St�$�3���~�@	�'��S`�̥3��\����
�9	�'@�i��WV7���b@�35��'���C�@�+��	�:������ Xؘ��G�	���٤ʀc"�Z"O9�4j�#��!X
ǳQ����p�O������́W|n$����rŢ��������?��xs�H��}��8%,ï�!�dG�;�)�@"�%o�`(��*F�!��h	�<����{c��KDMc�!�D�N̺YW��;#Q�ʓ)�u�J�l�_����"N�(Gf����/(����0�y��wɨH��)ޫ&��t������'9ў�(��6i=s���#݅k��ە"O<P�2H���h�câ	�,(�"O�y���4a���b��)���#b"O���֙6�9�g)�OĔ��v�i�𤍏=*` �����X��@
X!��Q���b$�ܘ�\�g�=K!��ً)��8�*�.6��L�1��Ą�t�ؽ��ȝ�:Y�1f�2ti@C�	�(t�Z�"�5��ԃ^�hmDz��ꒊه2���f�O(2ޘ	���1D�P;P�Ҙ2��))Ӥ�_\�M�C�Of��hO�����g�(�
5�'�X=����'��I4%J����ץB���[w눗a&C�ɦD���9e�\�_z�u����>r�\#<�r�'�?��PC��h�@a��Բ$3��!�@4D���J��%�� E�ބ<�����O��=���HOfM5��RM��8��UJ�
�"O.�pZ(�ђnB��9�w�*+!�dV??�䠠�ߛe�Ba��(P9a|R�|��6P��W�L�P*S'�9�'E�{r�5$�^e����7.�B��R����x�'��0Ń�s�-�1HҀ�jء�'�\�6 �&/�B��$�I�I�'0��� _�|ͻV�Ρ�P�
�'ߚi���g���y���b���O�����$8>���딶E� �P�ާlTa{�R����:ǰ�����4����b��ai3D�x0�J 2O���H�/X\�R��-��hO�OBՠ!���zA�Dm&4�B�	?*�Т�_p�.m��d*KA�B�I�ItE��˺ \F�˕n�B��72��=`���{xe��h�&J�C�	$U ����F ��csI%I&���z?IJ>"`�5.�\�;6��.v�܀1�s�<����F9�3T�J)C�8��Hl�d"�S�'8dpؔB[�jHL��
5b�܅�xa��h妙5D=��)")\0M2�Ņ�RF�kFAؾW*L����H�ȓi��U`�K(x^T�a��$%A��s�m��WC�}*g��+
$фȓ@	b5�g��d�Ԝ�E!�]D��	����Ҁ	E���I��h�ԇ���Xs���`d��T�L�j�̭�ȓ7WD��a �;+�r�Cn�z�:��ȓN�J��"���A& y�(���r�d�Ia �,	wƩ)�ܾZ�d���y��᳃živ��9v�
�O)�Մ�ZdV�	��@1��L31M�8� %�ȓT5�ph�O�0~Z��D�TR'�)�ȓI��1�	`��C&ͬh��|��As�d��
͵Vf�x
S�ނi� h����SÅ�-P���v��3l�� �ȓU��s#a�'VI�kZQ���T"OƑb#��0<W&�0�%E;K����"On4��h��$�@C������!"O� �����/gjv��e$C�Zp��"O^�1�o^:d|��B��r�x�Yf"O^�[�+3�ՊЮ����c�"O���ff�4{�(�1�S<���"OF��#Ѧ8�~�@ O�f J�b"O4�(�I/n :���7C��D��"O�ȃ�pN�	r�L�8,�IPU"OJ��O�%ĜHR��۵k�����"O)�4l�5Q�"�S L��b��4{�"O�]����L@������u=�Y�""O�U�Η�2�f�@49'T� t"O��s��F��i���1���V"OhT�p̜>"�9����%�l��"O�h�ʞ&I
,`��ҁ/ൡ�"Ob���,]�E%0�%�V5�d�D"O�I���E� �!�;~��pS�"O�h��b���|���}����"O���#N>���(��W�
�R"O�h�a��_����1�U ��)��"O09�p�'F�ܸ�甐L9X�e"O��Aҋ�>�΄��ȶC&l��"O )���Gf
�g�ȽOp���"O�����ۺ�ܜB�ő�ir�%��"O�0�cM����cn�52,��q"Ol��$��Skl��V�Y��r6"O*`8�*?]Nd$�A��p��"O�����.���6�1�><9"O isuD׼G��r��!�J0�"OR ��m8�F��@�Үk�$��"OJ�����,?d~@lōEJ���"Of�9�윇Q�p-�!��=(�DE[�"OfX2�i̚�-���	��x@"O�@�7oϸ~ޜ��h˱J�dqJT"OtY�ǓO F,�T�����p�"O�0{F��+�He�m�X�8�	�"O����'�6N �%��˓�w�P30"O�����A#B��5��& �&e!t"O@
�GQRL���/	�n��t��"OB�k�hN�:rF��m�:r���ٲ"O�h�`��9���� b�vTH�"O�d���훷K�F��a��"ON�I3�ؠ��� p���� "O�Q��\�}7*�S�M�+����"O�]Yl	:d\=ڱ��8���U"O���L�U�zwnE�2v���"O6!�b�.#6��ZU�Q
p6P�"O�qP�Hƪ#,����F�w�Bm��"O�pi��Y,-��P���}� L�v���<�!I�=-�N�����%����$Qp�<y��b���y���J(�[��Jm쓷hO�O}�`�U�䊣u� Br6era�4D��1�q`���#$@ p�j�O&�D�r���OM\l(�b�5-Pݫ@��9Ԫ ��'
XLPBD4��<����:������+<O.|�wj+{��� S,@V�YSf�'|qOU�'�� �P���A	u���H&"OV	����
�Y�b�9۰
�9O���$M 7�ȹ���ݿQ�,�jTMF�?�!�$Ģq��Y�� ިB�l� dL��ly!�D#ER�Ȣ6��3<�N´L\�x@!�Ě�R��&�"{�у˅�?!�Ӵa��LZ��( 
��J�!�N�}@�Ě�K�\�e:�	Ȫ�!�$�dd|�Q@��h�@�
.�O ���?� �����B�2��p��΂��8�*��'��qmZ`e�}u*�1$��BE��~Px�O�=�}�u�^�a/ ��芚u+P�2���H�<	C1<���� %ד��b��O�<���O�R��XY�N0F�0q�FH<qL�)3:�8�"�+�y"?J��HʣQ�h$����'�̝����B�V9h5� 6X���3�'1O���|B��DI 	T�|:eF1N�h��ÄB��p=��}��!4Xf��K&K����`��%@��Dx��b��'2(�O�,`�JX�l�p���GD��IT"O��f�1�T�e�Md�HV"O�I��>:JRI�#��95:�Q��o���)���h�B4�=M����ϯ'�!�d��YY(]���Z�#<�(�
����'m����Zz��G�\#6�R �f.�|�x�@��M���7�@�B�K?��Of�ȋ���
;�]�a؏�,�E�ͅ�Q��E{*�����L$�,�1������#"O�X�P.M,=��$ΜT�����' 1O��d�}����-"+$�QrC�6 !�ėv�̕�4��QL(�	��x� c�8I�ҎC1W��3�]�vX�m{�'5�܈��ʊfT�ۧ�V(t��1q�':�6�)ڧ|� ����9���[2.�@�\F|r��g�N)QF��a��|w�ʎf�ĒO����E!K L+'m��il&YJ'n�j5!��I�^Y��$&�W��E�cq�	�'.�����
Ih���/e��Q��hORY0G��J�
�X��FB��$X"OX(�0��lҌZ%jѠ/Y��XX��l�b��(�r��3�����BќwT��ӧ"O&t�ĉ*H>�!{�ѯx9��՟|��Q��F{ʟt�Q�n�n�  K��x44�9��'��>V7��CŀJ�4m��A�.�B�ɲ�x�qBҸ)L �J��D�C�t�����EK�.K���eg/О��d��$ٳJPI�8K��M�����1b#D�l�b�_A6�X��E0'\f�C=�Ѩ�<,�sa�mj�"��fH1��O��I]�D<�&T�u�p,�,.�D�Y5��k������"v��;'X(��'����n�A�����6��Ej6�A�	�)���`!
��?��'&^|2�`2��Y4�JY���<��D!�OΡ��`�\v=3��)t^�¡�I�MJ?�8������р�o��ٓB.D�$9�Hެ~��؁�CE�w�̘�$2��hO�-D\�$��2� г���U���>��`.�'s�������}f�-�'R��z���`�@�#��0J���{%�Q�%.:��I7R��?�'�O�|R%0!{�Ģ&���,H�q��'��IL~RMP�E�X���Ǔ�8 r"[
�䓸hO�2�D/8�%�#��J�m�6���'����)�Ӧx�>�5B �w)�X  �΋ra&lr��.��"~���uR�`3t�&r�q��˿k��C䉣�؀#��H<A�[ԠI
o��C�ɾ���S��eN��ۗ��˓�0?���� ��u�|f���/�qyB�'A�ɓI1z!"�C�L�|�2�e?C��e����Ѡ�>}|4k�cE:l�B��%���D@�(d���%��Us��PG{J~b��r?Z<�C$ݤ]��m�q�_`�<I�O�_��
6BƤ$~4Ȓ�D�<��#M�i3�F�U����Vi}��'��DGj���:A���1�$Qu�\���8O,c�� ��#���5��Yp���v"!�V��
1��'+�'$�}�Q��t�h(wM0���p�'��O�9�4���떻"�&5bo�f�V����0�'�V�Opq�l��k� a�b�>~�.�KE�'-��I�k�*1Cu��U�^�I��,�B�	I9��ñbш10t�0�)` ���>���܀@ؘ %�>74�pc���=�0>yq�8?�sb�6Q66���k�L�\�03I�u�<�ԃ�Qo�Z�9k����"!�[�'%��E�T+(#w��Ц�h�L��Ӡ���y"e��&_��	FYׂ} ��*�yB�D�������G�]��K!U1�y���gݐ����
\�p�����y�'8c�t��5�1U���EP5�y�ޓ�}ye�βMi.h��y�dR.]���E'�0��A@7�y�M�n�f�8&�N�D�)��$���yR�ۈR�Neaeb��pU�-�D���y"�90�
Y �N�8XF1P�����y��Yf8�
�9A.��� M�y�#υU,,��V��6�H��h�!�yҫі0�Z�9A`�-��,��G��yB�]<&�
A@V�+�l�e#�8�y�F�4t��SwM7y�<�E��y���|`qA�Ԕvm���T�ӹ�y�ާ���l��k�Ѕ���V�y"��t�d��O�-]M�5�R�*�y)A�y�b��7�?s�����V��y�a�Y�
t��"�.�j�)�B�1�y�Ğ�!�\��&����l�Ad��y2��79���.M�^f\���ݎ�y��͒�z�Pć��Kb�(�Q��yB�sB�%�teĹJ��� ��ʽ��IPX�x�P�X��乺2�D�
d;6�#D��u�8I���iB��
=y��-D�|�wl�i��Y�E�ۧS��yjs	̧T��7�)�矈j׆#,T��Q��7��0&-4���4��C�4��-���i��J[A?q�'n�YY  ;M��k��8���r���4��:�`H�9eH�n�	q�C�I?��p�pnѦ& h
TȈ2y�B�I�;��%�oK^��a)�`��Z9�B�	�cK,<��d�1�ډC�L��7�B䉭!����R�~Uh̹���7�nB�ɁvIj��� Q0O�*h��눬uh��ƓYev�Q��!2J���(CV��ȓ'=��*Rˇ)������P��ć�U����ď�zh|[s"Z�Yd�p�ȓ$[��`�C@&'����B����ȓIu��X�n����uSu�L�!`�0�ȓ1 .���ě�&U۰L��Y�ȄȓD�b�[�,I�����W*%��ȓ^Qj��C��F^r���
w6>�ȓla,�#¥��l���s��VZ<f�ȓ��ۂk�>��5��g��l���ȓ2)̀����dT�aʆ,��ȓM����B�@�RF���7G �����w"8���7H$���A�:��ȓD��<�K�"j	�1鏸DL����X��O�%)B�v�&1~y�ȓMRu�r�*:���ݳEi�E��a�`�P��a�dt��M�dގ���V�&=��l[�+S~ �b��=C�Ұ�ȓ �d���ϡD>��j98���S�? D,�7�K���@Yu����"O�x��ϒe ���`�*=�X@@�"Ox9ˢz������&X�4:"O"| 
`8Za*u���$"O<�� NH,�|57"�+�bdS�"O(��I�X�����.Z�gTth�V"O�����'��C�-rK4�8�"O���@Q��>��0↛|��i	�"O<�Aԧ�k��dSt�D����"O�,��FC� ����q�ҋi��qc"O��h`�I4q���2B�F>�1{�'��4[�k��'����m�e̐�r�'���w _ 2t��S�U�W'̔��'���ҴnZ�/�x�Ã�ŦS��p
�'���v,Ӥ.�d�!nH6Lh�@�	�'�lE�2.^���` O�rg
���'T�l�lŰV R�jK�l�����'�����/0\�j�Ń�{�L��'�ʔcU*>�$�{$��+�,	�'�~e� ���f�p��A���0��'���"7�'E� 
ĮI1�ڈ�	�'X�	s���f�� 4�ݢ��l��`7��&��E��{©O )��$:����Ok�B��N4�y��F �Ny(�-@=G�n�B,�y���?ɒ 8Si�:Ԣݚ���y2+M?M|<@�e�2b��hE��y�4��@a������ 2�yR@�=�b�@���$S���ybQ�8��Q��S*���h��y� G�f������:Ag�����y�ܠa�n�ö��V3"��a)���yүV�2��yٕ�L�VHQ�+�+�y��&%���K�9^�U0� 9�y�سh�Yy򣃲?�(�a ��yr���r�&��Q��/�(�raF�y� P�*i|%�	�%�&��v�
�y��
.G�Ф"�,�`��5�P��y��ʘ�b���<Hؐ����|�C��+6頥`�^!&0�TJF�\�"C�I	(㐹�P���k�@��=M(C�I*~��4f�G�k���g�-a� C�	�W��A+NI!}r�#7��nA8C�ɞ`g��[ۥ]��}��O&8?��K�A����S�O^(00������.:j0(R�"OXL$�?�
= aa�pVȁyAŅD��B�!妄+�*����@+~ �^x8XYCE!da2��2/�Xܘ�P&��\��}_� 1I
��q��'�ll�lѮA��!��L/I18��$��f�b%*7O�:Va~�O ��:$�|���K���#C|��2�'.����
���!�Ì�v5��X�ODD�Ŧ�j��1��z>9�g�5}P !'%����!�1D�T���of�5f�/b�~��w���j�����7	��L�9���%>�yҷ�r�	#_d����P�9/za�叞2�"�� ����hghˀY�T{��]b\���	�w�� �E��5�<��s���"�i&���M�k�'���s�g�,ߨP[iƟo�VA�7*K$9�H� /��E�l8��'K~��IR�#(�$��<����G�8���C�I�>�1D�8��	�Ϟ�M�\#*C�D���*�	0U � b�I � y��Ա0�!���p�b$��k *&��e�'��A!��Ɠ;��aЂ<\(X���"=_ʓ�r��rl��o�b鱰���G������v���9w\n��+0E�$� 5B**�ޘc�e� ;��!TK�Q&L����I�\.�&M(���堅�S�����[VDy�+юY>��5���wy2�K&ͅ�d�����^���k��<����/\¬�W�){~9�>�Sꁟ\I�
�L�6n�l9��ߡ��3� t<zfC�ptkP×�M��d�Dӹ;[����9�'1P<t��.�g#�h#@@}�~T0SC{����
2
 ���E�O>����9�|��w�A82&�QF�ٓxR���l)��'�4�|�'�(2�B��)��;E��)��������.���b�O3_����h�8�u��ɯVu�p�u��H=��n��[���z'̶_�����ΔC�'�J)��n%^����G��"��̃�gn(=�tIF�N'�uP��ª0�Q� X��S!M�pL���ǟ���'�U�,����-�Vd��9�I>݈%3BB	*d����԰䧟n ¦�H�'N�	�o������$���ȋj��o���}��S<����K'�@)��O&T45��(��̸�I�P���}��'&XB�Ɣ7�4�	��ʱ+�ԫ�bD�SbXeۇ^�8�#�3�g~����NL1�l��@��f��E�� 0HdY
&
ωc��D�q���3�{�F��0`�W5!A91`M�.$T�`���=?�vIC�d��p�:`�I��p(���g���&��g?���O�v��Y����m4�b���I6�%��e zxҝ�&�I	��d�Im�)�n�&W��q7�G�����@� ��d#�N�LS��t���j�(���Q:3�)�݂�M�w���{_)rf �5#��c 
Ď{נ�|��X�P��N*I���7�
�~��݂��<⨘�D�yw����S��y�i
��x�7��B���`�[����3�
��U��{�˟���먟��GxGM�El��U�$P�#���*p��V
_��cB�Ż�x��g͖Dl���Oڑ@fk̖>f�:+S���E"��
J�h��&�4`�6}kA��$�"?IT��8�����-n �<h熇<
X&,��#@>ش���wjr܋�%�b?���i�c�^��O�r(ks�D?h�`#*]}�ٍ�D���2�O���O��	؄&��I����g��h�� ��4 �ތ�0~���q@���<�'I���㷇C�$�9+E!y��ƇC侘�F+�N{�$�+M6<*�{J|�UDG�8;�yB���Z�v9I��B�A�-��%�6`�	�&(>�K$�P0/_z��	�9V
���,�
�Ek&0m��=�R��D�b�XAk�Ԋ�Ɍ+7�D�E���i�:N�N�� X����'\lDz���"���b��to�-(��F*�A@�ۭu�d�	/2()R�C�q���T�6Ǡm��L�d�n�Kqi>D��
3lم4�i�5Gǚ0�&-k�f�X�`_�X{h�ic������O����c�,�DmZ����0Df5@'K�n3�}"�ˢj9 �����A!ٱ'�Ə}�Uҍ��
`��/��ɁĆ��;8�P1D&N�^�G{�<nu.�Q4�NN�(�N�3kٸi��L�GL �>�Ľ�ȓ�H*� ��R^쉄�P
~��y�2
:| e`E�~���\�7m�S\���
��q���r�΁���UJ¤�f��Gar��
�b�@c[:EaJ%Q$��wd� o֑
1��CDF��F�� ��h�P�O`N-AK�C�]?8G�]��HT76Ql�Rp"�Z&�C�*�52���"ER��V	ܩG =��٢+�i2��h�΁�!Dp>1"�b�!BqO�0j�lH�"  i!o�C�v��g�'� ��]<wS+��H}̬�e�H9h@��E�i<��L�uS�����T��Pp�c��Z��-A��G!@�#;a��I� �F��2;"B׎/G�Dk����	p�S��E�5j|�S�W�&	����,�p�<�WN�B{:����Ŧ�S�%� ���ѓ�NY���+��Z��Y0O�=��|�}�;=�a�Fa;~�ؑ*!G��?�|��s�fm c�\�)H��G҆
�j�#7�V7�܅�$Qnu<]ȐJ��|3Mܺ/D㞜ಫ��]���b���HFE�j;�OU��j��R�BP�u%�dO �CgI�L-�|h� q���y�Dб>|�\�T̆�p=���E�Ne�|�4�3W�jzfDR�'Έ�pr��7������2g���8�,H'�ԹH�Pޤ��D��O߲�c�(�y@q]��@2��k>��'����$8�EH&Qĵ��#�8p�!@�Ls_��>�;� ��A̅o ;B��3Y���zU�E�rJ�2�a �̄�ͪweY+��AA��R��D( ��K6�J�>AR��$D�)O�8�Z�oCu<�� �9lO�}�"�;�)��))x�qr�m�t<h ʕ����&�P�&�C�(P�'�'D�8l�M_=[3�3�6�I�s�Լ�e *�M�-�4|�`�(GȌ�[����(|(ډI���Z����
��y⫃>>�������5]�X3�hV([�.؛[��s榚/x��	S�+U.Z�ᱏ�4jvޕJ�iL2K Z��d뒢�4m)�h9D��[�-� �ŁeCW�N�X�F�T�@��<���]1~��dKŐlsD�]66�p��֕g����u�ײP�,�JT�SDMa{2J$V�>X
�I�)ɦ���D�<.僣�9`��!A��F.+F�p@S==����t�,a��]Cx��ަ
z�b����iB/��U� D�	Tn=�5.O/~�>���Oތ`��L%�E��P���s�\O�<�ō�6�{�E�R�4i��_�R���CиBy.�8��D�J����EM���O+�� 8�piU�z����+�/%�P���"O��r�ń�`S  �׫ͽ�fp�h�t^@�3Fł x���#p��X����aV.�h��/����Ԫ��*���V-bӢ�e�Z��X�?A��ݷl,Q��H�%(yZ( �M!a�����pu�g��"=���	 a����Q+�	�Ĉ,����p�A+#H����(8�����I�be�@Հ!@u�
T\�0
��`�� "����V@̓"���j���j�)��)ك$�E³�U����DM�I���d�Lr���`C�AV����������I�U��<��Lc�P8V�-��l
�M2z{��!>Y�"|�'q��T,�'E�(Y���3Z���.�~�	�?I��X��V� zr�Ef]^��t�Q�DQ����K5Hb�y���H���h4�	�$Z�U:���-a:İy`��
x"���vm?=	�鉼b�D��폜���� �8EcB�FKl����̣@T">�4$��iNj�|�v��A�]���;#�X��H�j�&�p�Ȗ�k� �Ј�i�9Zv\������>�D�&\�3�1O@�6$<<O�,���da�T��+T�)U6`�'O d��qVf�<���\����	�5���WgŐ4�(@ ��(�!�D���܀�ԩ�=ZA�LR&h60��*�O������5|O.�`4o���B�7bP�;!�'���˱-��V�JL͓6�<�h��X;K� H����Z�d��\`Lh�F�(���`�͑�u�>IS���B�t�9���ˌP��SPdݩo �]��"аd�!��A	Yp��Ap�`Rt��_�L�!�F�i���ƀ`Z� �Ήh�!�DY� �����.�٩�S�9a!�DP�rW@�:�L�Xp ���g��GX!��T$��|Ym�$I*�c �O�INAF{���'�bUkR'FL@a�r _�z��|�	�'�����Ϸe5�Q�R��M��0�'a�牴f?��%GO1IE�@�����p>yJ<i�C�<�\�HQk��^ӤX�C�NI�<I��ٹn�K �@"7�L��i�E�'�ў�'.�V�B %-m\���mϽ�!���1���I�@�vg��9C� ��E{���' RD���v��y�R�Y���[�'< �r��v�r)!s ��Y8���'�a�ٴ=��Ҭ�=q*�Eb4�p>�H<�rhPh�C��^U
a�!�Sg�<�Q_�f嚠{��\%4*CCV�<9��/z�hq�p�F~�Ұ��$(D��A� #s1�  �@ �dH���6�%D�����6�R�P�@�W����i6D��� *�%
����
�Q>`��F�3D���BѪ ���Q��)�Hp�/D��1�[�D�����h�O&8��m>D�(�6�@�\�J��j�9?{lx�t�(D��V$�<>��*"a̺}0�cg�0D� �5l�����1�,� ,]��o;D���P��xM�ԊȪ2J�Ѷ;D��BjRxT:M!F��A��dD,D�D��JGK�`�Ǥ5ުUR�-D��1��\,�����I�& ��Cn,D��b�,6k��\2q���FWny���-D���ѣ���>��Xq�Te9�l�8�y�aO*u �T��GK+~���F��yK<#��R����R�0�l�:�y�F�=j�$��zN����)]��y���1$��h#�j[=rK��%�ŕ�y��4&&mk`U jt$���E��y��:�R=@6f�l�Ν�th&�yrjL|(&�Y6�vh�����˞�yA,,��m(����ӭĈ�y2����E3+483f
,/!��6mV$�2�L�r8.YO���'u� *t�<=;�8�$�M1��
��� ��)k��Ӛ�+¬��Jt.�4"O��A��Q�#g��K��Ȅ@dZ��"O �`a��z��ⳋ 4l�D"O���NR"km�A�"��Z�Ę�"OB�U5���$�$xN��"O`P�j�J�Gm
�M���@�"O�]ke�B0Z�� E�
 �dJ"O6`d�_;M
��t�L�!��"O���]�Mi7i�X�c�߽�!��Æ�֭yb�̊c�`|i�o�?t�!�D	����+B=9`� `��)�!��>~\p�˖�0R����M�!��U�m��x��'B��lڲ���v�!�d
%CiqRX:�(\�� ��@!!��H>_e������.S��T��J٧S�!���7#d3Θ8A�\��P��!�!�΂YF p��@P!B�1�Bf��!�D�
dF�شg��':��;TE��g�!�d��	G���7&�)�e��o!��,WHT���	&��03p!��,q;�=�@��W x
�$��!�ĉ/p��
r*�Z������@�!�D+�4c�̅4f���A�!�DV�^/D���,[q�>�Ac!-2}!�ĕE�x9��Ҷ#��|�B�-jG!���B|h��/]x�
��a�c!�$��Q�
a�7�͙�|�[�`Y5G�!�Ď�;]��1A��N5�ċ��N�!�D��3�,%���2��e�&���!򄏶=%�#b�GCe  8��W�!�dP�
9���hD�t���Rj�!�d��0�I8�`ƅ�$51���f!�DL�i���@B�ۼW��a��N�!�d�"	�t���M2U[�]8�QJ�!���&2��(�����N[ �@Vb٬s�!��И�C�@ř7@Hx fk	�|!�DR�r#`��զڌ[4ҽ UɝPZ!�U<$Q���"�M�'?� ©��7K!�DN�l�v-g�������\5!�$�-o��jt(U�d���2��k!���V����IZ^��ځK�1!��]&ͱvÛ�y0�-H�*��t!�$�q��$�afϬ7ׂ��Љ�e!�}���`%ËuQ�0�E(� FN!򤐮���i��k��2�i8�!��=x�	�3�K^F,E�Gk!�$R@���T#�Z�����爐��	4��UQ��Q�)�'��|Y�b�a��5�Qi�j%Jчȓo'��w��k��$�󫄗/oBm�f�>Avg�-ZԐ�N~�=��E��T���k��6{BŀtAAm؟,��K�"ͤɢ������6ǐ�U�A���Z-yTx���	�H!Ӷ�
.�:�:OEy}N#?�ʙ�\d��T	՘����Y�(+G�ԥE��x�g�=H4.C�ɺD����R�)Kb�@�i
)j�6�Kcv`9ңIYFE���O3�1 �I�la�4�Q�'?0 @�'��4Ri�\�]�QF���K�SyR�̹'Hzta�+���.C��<9f'Eq� �1�+1`=a"GY�X%K*�7^��t�$L-qxU��EV�2��d�5�'��@��i }��Y�B�J�Ix8c��D��M��;���S��O�Bm�soT�M�Ԡ���O	I����
�'|���R��ر���f��O�t�v N�����W>��"��!�T�sc]��B It�"D������;h(�!rdTr�Uq�+C�����	���WG�3�	:oPQ�Vc�-+�@����аj�B�I:n
T� �����I�*C���G��8aqϽ.�����K~p5���3<O>�ꒉK4r����ը�x'�M+��'&�]�C�-,��=`��1c:����S:��Z�m�CH<1rd��f3f��05+�px�j�'dT	�,�24��`��i��UD��Rq/l\�H�����O쓁,���T�~�t�[�&��+��a�^禕�Py_*�Q[.��S��M��*I�[�z% g��}�(��_"������B���(��Iu���pg�i���Eb���3�O���e��<C!�8S�<O���I^��\3P/�	E� �@��b���C AL�� �>AD��k��@vI��m �듌�9>�@)���ݙOl���	�/��HS�סro2�9��^�I�3g���u)�G2yEz��\Q��E�ƒ����a�,'��9��NB!�Q����ט'#�R`��Q�Z"�k|#���Ӽ)�r�˟q�\7-��l,B��#�5FW*�S��M+�n�u;��f!�1c9��2�����^�;�ȁ����>�)�0Q��cy�-�E���r�˺>9�a؟y�h��	3�(O�9��
:Np܁w��ݖ�����+�.`sJ��{-B�!툞o��#?)T��R?��K���8=�� ��]���&�&_~�<	�e��?��#�l���-�<���'d3>D8�-J [
�8�B�PL%G|�,F�	��Mp���*�"���	_�6��0�ĭɛVE�3^6�� �������ٖQAF�\c����QkT�k�u���	mL��2�'�~(�T�ԧ*����iЃ_ *��`OǃM�F}��O[*��e R����ST�'J��Y�J�g�� gN�H�� C��̞$��y�O�T�u�#m�!Q傖nW8��E������+��P*`�V�^�����܂[� 	��Pdib��$�^��a���p� .�.x�բ7��r�'>�*�󨞧v��@�7�;*��p��:���iSۊ3q���M7'�R�lZ�1j>P3��Q~����${����2t��c�-}��ТT����vJP4иpAs�ˇ��>Q3'˅�z%���T���11��9c���#��9�.�	5��c�*�<6 ����
R�� b
��J�f5����+�6�=��b7<���1�r� s3'
-N,FEc����Q��.Tl�5˽�D��(��K��.0�.��A��^��p��86���z��C*f����ȱ)�¸O�~����N�cò�C�̄�t`��"O�I`Ђ�;K<�*gJֳ:�
)�0OJ���$��v�~���Q}��$�@�S�|�Z,ae�����g�v�T�>��>���<uz��"��I>��%�@��[[���cn�w˘B�ɵt�F�s&�XviA�&�Dad�=�Q��4R�ҝ!$	6�ӏi��0��̦�B5�EKO,I]FB�>xBak�Q�p��B��J5}�I�'�!wa�h?� ������ѝq����4���;f�8c�A5:�"����J���B䉗C��T3�ɞ�-��u���nx1���1���"L8�?a�n�A��\;�'-��U�?��7~������[�a�J "{-!�����'P���@�bR�38��Z�f�h�+/,�@��y��)M�R���x�{r��L��e��%S���	� ��0>�5�N� �HD��$4~�y�ChD3:���5L۶q:��c��;�Jt`#�\ǰ��dʇo���PO֭S�R)��c����D���ܗ	�n%!��^��z"��;!�Q�Э�?����&J���:��'�Ûx\`C�I*Q�|���m��t��]0g�ͫ1z�:U��<i�b�g��v�д2�P�V�h����9��}��vne�'*Y-@�1I�"Oցx1��e��5��J�@[�H6)]	Y�i6I����ht% g�󩙅f���{B�\r[����;8.,◣�8�0>�1��ұ�V��Ua�m�(k��t�ǫ�2j�`�8%�\ܚ��VON%~������=eO��I&�RA�ְ	2�G�AV��e�6x͒��㬜�/�2�qC��Y��d���	"2u:!S��L!q)Q� Q�)��B�& kr���痯]4ư2c��9|Ba"���M{v���L*14�ܘ�ԧnz����:� pX�B�p��p��̥���q"O�xfC��=
&P�6���n�t�4*
�a6����nQڠ��`ȧO��.�+��4��B ͽE
%	7��t5�9��'��=��n�8͂��d��O6�򱡛�4x��F��}�
 ��'�9c�g0m�a|��2$�Z�q�k˕w�(V�ل��'(�	(��_�̚tk�ɮ,U^�	�B��d���,5j%beK[=%P�"U��0B�I�n�FhQf��!Wy��QPR`�ب�担`�z��^�@(�A�k̹j�N`�}��6����ǫ1 �X��n�"��Ҡ"O����!��X�3��jb�Q�"�	Muz H��	'?�~$�FF�$/D�bp�)�I�_<ܡӁ%]�n�J`CK�\���M6Cx@9�C�
|�t�� �Ш���+J�$�7��6E�a&��/��a�R�ː}&���.A�%qN�>^)"�F_�O
�
db�O�R���D;;�D@Q+D*i��'�%�C� 6:�ID�pd���&�l$��kIDX���p͋�K��dpBiJ���e�ؤ ��ˍ#�`4����1���u!_l�����6;$���"OLP�3��a���A�T/a�mC�+��?�2P#�	�xP�*VA�5b��Ƀ�`���(d�Z�^�r�G6l�|1�p�n0rc�X�]l�?�K�n��)�A��Z,"���CzU� *+6Xbl*&��<z��&�M�'3�8P�R�4\fhΓIE�d1E�ߜ$n`0
��_�p�Ez�H�'V��򠯎�47c�o�9��I6ئ@x�nQ
Ъ�=x�1OlY"�JN�{�j�H3 1ڧ��d�u����"������kV�hoZ�.���╠�p~ �U�j�"~nڶ�J�:�./�6`�@��?c<Ek酯'���'D�����Bb��<���Y	 � )pda?��MKh�'�ȁ"�
�?1eL�
Q�AAK	!��r�,R�J���ER�����#l�j�:v*D�.��S�K�9D2F!QER&��d��!�%�`��*�v�dǏbo����!G+��m�vf:����q��_�Q>��rf�2_P4�� 	�q�80��2�8sx�PT/�9,` G��BR�{K211��k�Ʃ9���"�y����m��t!0͔�
�'��vQN!�F)� ��	0�#|�O"q��O)V�
 ��#hl
���' ��5O3EƠ2'�ơu�6�)�΁[�z-�!�L+rC�{"۹XY��▊o��p�M�p=��b��j;�i�#'n���U�ݧh�8R�)Y>��n#D�(s��TlzN8� eE�xU�7�,��2_��*��Eb�O�2����٢9|%�q/R'H����	�'��MɄ�ş1Ŧ����\�|F�J	�'�e��
J��%Ò+O� @��'8>�X��c}v]��*��qS�'d�]�.��$PFDI�Q�ҽ��'������5U�d� ��H�?u Т�'FȔ#��?*�F�D��$\V�Q�'kHU�cEҝ.@��C�g(+G<A�'K�\C�Y#7" x��lϯ%oV@�'��b�Y!/��K��N?�����'Q�`a�LR�1#��j�v��'�4�s�Fށa�@e�傎1x�PA�'��Yq�h��Zآ�ͅ�xBj�!�'��lc���XI���bƤ$}��'x��D�J�l�;�aɕ(Y
���'��Z�e�V&G?+Rb��b-Ҭ�yb�=�dBB�#���q����y҈?yԈ�R�R�{���cB��y2�O�V��)	���:4�IC��=�y���iH:<$$�%,�d
�B��y��<d�����Eu��s���y�cL/1aD�X�À>_�2vN��y/�'&��,p�Û-E�4��ӷ�yrEO��N�P ����d��y㕵G�*t����3�` UA�`�<��]�[A������D�<i�$�-U:�U��@@�mB&Q[��
G�<���R#�]�R*ոT���4À_�<)��Y%�z�x�nF6T��pc�X�<��M(�&��2`#:<�r��U�<�a�,%6�1R��.Q��h��#�P�<)V�J]����+!r�8f'H�<�w��6��(��ί
���s�FO�<сD݉w�B��#�cd2C@n�<i�c��1φecW�ӱb������}�<iN�5�:PrR��eˈY�"�G�<1"h�k2>lI1��?4��#g}�<�N�_���cm�'�V�0��[t�<�e�/L=�v�9���0��x�<����oB&pb�N�_@���R�<� B��V�/؄�b�k�9�\i�"O���Q��7�����	n4�q"OL�D�U�r,z5�,Y8��"OBT�+�	�R(AFCy'6�ك"O���T�(����E�D.w��Ҵ"O�p+F�J����qnňx>��r"O6`�� @�jpX4^���6"O��9�?s��ʓ$F�v\����"O�(��E�=���Ѳ��#,gF1Q�"Ojq�ű3B�� fBd�"O�ͺ��ط5��DgC��'kr�A�"O�\ p��({�����\V Q��"OVuI֢M	C|������?p!L��"O�e���4| ��fS�QH��Q"O8e�G7i�F� ���tQ�5@�"O��yeN��Ubǭ<*XZ԰C"O�C���.0V̙�DJ.�ˠ"OH� 4b�����J�7IL����"O88�V�W���j0�w.d� "O�e��/��7�~pH�jϙm��4� "O>U0e�ߚ,~�Y'���tE�s"Oha��vzص��k�"��P�"O��%@�7-Yڥ§+�;J�@�1"O6�q�S2V���Diӭ
t�$x�"O^��0恗W<��!�g�Ր�"O~9+��D(�� bsa�+@а�P"O��I�3/� ��ג��53S"OT3r�}_d��UN������G"O�"t��<����$�;�4�3"O�
�3GD(�l������A�ߜ ����E�
�'.�=	hI��&?Y��%9H���i�
�\%���%8X����Xa�d�>��c��"c$���L�4n��	��9�)�?���P�N�p�L.]z�m	V	�@���?��\��y�O�(�(GL�;��
�ȃ2�&�8��$>�S�$	�,����+A�S�`I���3��'R�I|>�5���'ϲ�BQ	t6�qU&??��O
b��'��ת8H�`%�E�e4l���F�r���<ٰ-�>E�4M*�����$vB�[W�����$F���	�_G`I��B;l�T��c�6i^�����d��yB�}�R��c�M��p��E˰m�B�Ie��ݠa/ӟr�$�3Ш[�%j�C�	�X�D9�N��6[���a^�k`C�	sj�d�@��
 `�2��Z�`
�C�	������8��\I!���w�C�� ��1�C6��D T�@
c���INܓ�0|�F
i����'5f\R&l�<Q�I<�yb�ijD��Z6L�?�Cs��;k��� ���nb��Qu�c���`Gm�48�m�0��4����0��ħ{@�<��ǆ!{.�K�˽�虰���}}n�Ē?t��؃ш�I>��JD�@�p�,]���V��$�vLp5 V9n��@/l�H���O��A˱K8|�Ř "K�m:4��_4�V���Xxis��Ih�Lܧ|�Ji5�$j�Z��4]-ЀÇ>O,M���� �E��"Mx>]�d�P�5�P�д�\�o�D��Ê~ӎ���U���dě�y����4{�񖭓6���!AϿV�.I��@>�����=�)�$j��P�-҃���`��GdK���`��@Zay���M߬9ۅdӚW�ꈘ����y2���pܣq�A@}Vl*6�ɚ�y�@�)cb��Y�JM�>���b�d�)�y�ƞNhr�.Ӓ;L��!�ʽ�y"�D�<��"� ��=8D�\�yRK�' ax�LT	Ꜩ����y��<	H���A��RB�5g�Y$�Pyb"�..�`�̆�z��P%�g�<�Tl��q9rHS�mTz�MХ"M�<��G��h����
?�VX��Ec�<� :1��	M�J>p��Aƅ��0�"O��hV,'(�����*O��R�"O
���͈:����to��{0���"Op�:�¯~��z�g�	;�	�"O���ѹ$HИ ���p�&ճ�"O�L��/�	IU�܁rIFF��j�"O��qB�c��-��GA�I�f���"O�1;6�<(�$٪����N�� "O��i�OC<����d�� �h|9w"O�1q��"����ܻ�"���"Ob�W�̙R��D��T68g$�"�"O6�Y#��q����a�N,>�FI�3"O�U�p�F�9��1�Lߊ? b&"O�ӊՏB����R �P��"O�`��_l����	ފ��� T"O"��&��$��؂5�;3�4I�r"Oʍ���A�
=j��p3�M�d"O6�cv�L��Yq5�*b���p"O�[��	z��e�Ţ�0iW"OqA�~,���J�!����"O���SK�E�$��J
�*�6t�b"O,�*�D(S�T�)B*�e���Y7"O���b�Шy�)y7I�Bk^�ٵ"O��0� C�<�S���F�ԉ�"Op�B�Bq�,[���f̄��%"OPm�E���:r'B#i��USV�:�y�KL�J`a�̡gHr�rb B#�y��N \�`43�DH�^o"��4��y�bP.�(�g	C:(��bB#�y��q &QC�XE�x8d���y�"F<u,u(#��.����:�yB�R&e� }��O�"��q��+���y�hR�u��hrb�2��P-T�q��'`��Bd�-5��@���ˠ�	�'�XЁ�ȉ	:��1��͘�a��'&tؘT���8�}�A(M�A
�'Xu�4�$X<TJ��?;`|�	�'�X@���T}�y3�'��*�M�	�'LP9ЅG�Mi��B2Ϟ.TR�Qh�'�^�)��!~�d0���TX^=9�'�e�FO�����U0y~M�
�'䐤��Nb�2���Ɗ�4��'����4���A��S�q��1��'V�*A� +ypj�g�H�8�'>�%�Q�]�~3J(�������H�'� 1V��51l"�z K�\�q�'"������t��áB	���C�'^�%�G�գT���BaߋU�t���'�t����4_!�a�`@ƚ>rd�`�'�p�3�)6�I�O�b���"�"O���4�C%2�L ����3wfh�"O��b�*�*GԄP��(Ҕ_���"O������8)ˢY�@�ג]Y�J#"OX0 w�^j�Œ��ֹw�~a"Q"O^A��Ů�H�X�����uBw"OtM�&N����l
%#��W��c5"O$}�p�N�ԩ
�^=k��� "O��ȃJW%;S��E H�`Ҡ,*f"O�E�%��8`E��YE��$@f&H�#"O�MBReN>H�%��);R� �"O��c��Z97�1���˾r">L�"O����-Ģ&Z� �s�*4	��ZG"Ov�٧�[�t�@���L�^���h�"O.�����|�ޘjWG��>��1"O� �h�HH��.}0�'@�.�^���"OTi�_�'����� N�M{fU��"O�����Q6��`/3��ae"O�({��Z  ��/I�˘��"OR�%D;<;��al�\����"O������d��c����5����&"O�͸�iԃ4�-zv���x����"Op͹�,�E~��3L�;A��%��"O,m��B�*g8�`��"Ҽ�"O��r�'��D.�L&%P-$�t�D"O�5 �ݛew��n�9,> ��"O�ŀ�σm6�̭"\�j�H�M�V�<1�� as�5�".h|m�v��Q�<)�ON��`�Ye�*P��B1KP�<�/�>cT���	��s�@�G�<i�,P�l�
��V�F�Y���K�)	L�<)$���EWp�ؐkC�K𠔳2GS\�<W�¢q���1���<)���j�V�<Q��.V� P�RF�.d�nLb�&IP�<��.9�ؐ�/G������e�<!�$�4V��U��%؞O[$�B��\y�<	t@�,��!35�I�`Ȓ7�j�<�S�O�Z�&�� Q숕ʡęi�<��wҌ��#�@�gP����n�<ɥh�<0!�I4��5�n�P`�g�<!�e����ɶ�\��-"�ǔb�<���T�yt>Hs�lA0�9��^�<���6%��$KRD_���BZ�<i�$ D܈Fb�5	�AYp�F_�<9P�9�X%��t"*Uy�o�P�<9D��F ���ǈ^(����P�<��Nɬ ~��$	_�W�V�($�I�<qA�L�^�XA�e�J"�l�ȣ��D�<Y�O=rb�[㮎r��`�CJ�<1����&�
�ʆX^��I`�@F�<��-�02�Z�rT[�PP	� �<��D�
1���a��g�@��&T_�<Y5�Ѓ�,ڕNа4�z�8�*�A�<V�Z'���R�圡,�LQ��� t�<��m�b�n��#��J��)A�z�<yC�+I��b���1��O�<11%�-`s�@��E_2���@�I�<9F��-4�X�2��qpN0���_�<��+^ج(�+p�VIj@Y�<�p�34�R�f��2��iBS�<�0)'p<��j���h� #�V�<A��a��ׄ�5E�<��7(�F�<1v��[�Xy �#��R(*G�F�<Yc²��E���O�-�*�aC�F�<�CDT
M��D g�ц:Q�T���K�<!r�U,��j�f+�r�	w(l�<y��%D�@��"ţg
z)�B��h�<�paQ�F��I����.3�Lh��b�<���U9&�~��wo�#N4�j�C�<�Q�k0YA�ED%J*F-�j�C�<����{d�}hQ�� E5�T1��A�<)P��h��sd�6t��"H�<	T@U�!c�m�An�:wN�A!��N�<q@�t#R	���U/Og ���M�<	�#��s�&���qu:L���H�<I�LJ'^'���"B-*��2��A�<�B��+��\AR`C]���r��<�`��:`ᩆ��Y�f��*�}�<��EȲm�~� �S�6�j�mKz�<� z��vۮ&[���U�>A��Iiw"O��{�E� ��A֊�m��y�'"O���`���ji� �Ui�2S��)@"O"ݡRIۤS�+���9g+��j�"O^���Gҧ$�2�)�a�%r��"O�i�/� ��AA�����$"Oةq"�"X�2����7f���"O�]���2s
pe�f�/�\j�"On<YèJ�y#�%�� �� ���"O��*�e��P���eƏ�D�Q�s"O�Q��
��@���dĩW�4��"O��P 
�3*�d£#�^��L�5"O6X9���f��{���8S�1C�"ON����� �\�bT* ,Dpx�"O��0q*O��D�js6<qd"O0�����*��h0&Bl�L��d"O�Px`�R�Y��:p�L)h�p3"O��	'R�2j|��Ae܆*���"O��#�̓>jLiPs�ϕ *p�p�"O�(��΅I����B��;��Xu"ODIH4g�(4�@���(*�$��"O-�R
��~h����c�h��%"O�-q�(N�*�,p���T7�]��"O^H+���$��9���\.-Sh��3"O� �!d4��(s��kX�U��"O��!����\�ҍ�PV8B�1�b"OnЈ2晨Rʦ9A�@�;R��"O�,��+�:4�dL[`M��yq"Oby�de̤D|(���/�����"�"OJ��m��n|�0!��=z��q��"O���g�"���IfR�"Ox�B�,�+y�xd��3Sj��v"O�̂�K�t�	�������q"O���Kİy�T�����l)v"O����	TP�CR;1�xH� "O�l��G��YL��DB�z���+U"O�8k+FE~͓2/�~*��c"O�4��@q%� ��< �4Y!c"O��{A��W$�@A��07���"O0X��Ĥx��h�S/��Ҭ�"OF��`N-r�|2"�
����"O��Q�F�<0�h|�%&�.w��@�2"O���X�^��c���6R�ҹJ�"Oh�! 
"j���I,Or��&"O�a!uƕ�o�N�q2G�g_B4R�"OX���%�uQC��T�O�)s�"O\����>d��e)~@��6"O|]���4]ĉ�J)Z�F�Q"O�DHB#R&y�����(!!Ȭ��u"O� 2�R�I���s�|ءt"O\�s0ぴ��M��--"�4,@"OܙI$�
rp��[�fޛC�(8{�"O����U�,Ǭ0�6F����1K�"O��(2�d��iwb�0�J��7"O��j���Y.����@�m<���"O|lY�@�;S�)��	�Pc��ѣ"O�=����E�[�nϥ�@b*O�`��Ŕ)K*�=����.s�B���'�<<�q�94$�91�M�p�PT���۞<f*�oZ��n���M�'r�.� ��?A��MsY�<���A4�d�«G��,%a󈝏|{	��3Ҹd
S(�?Y�OW��@��<��"Iw�h��#�r�l�Е��IXq�'��mW|���g`���;�u�g%�iEļ7�ْ3>���fX,1��Y;p�"�'L�6-�O�=c��Y�(�+�e�^��P��%3v����^�?َR���&�ıj7� X�"�j��ڈ.5"�H�۴*2�����x6� \�2h��h��Q�2�\̲�����,�IR	"\N�I�h���D�ZwT�'���O�u���H1� K綔R�U�<m ���
 &�����1�iȓ!�"ψO��Qƒ�LƠ�AٟO�R	 �YKg��ڴ�S�x]�O[��Mc�/��a�D��}��+�p��E�4�y�Vo���Ms%c^ڟ,�I��ē�?����ēzrj����F�PlZL�0A®F�X��?i��?��H�`���)OX�d�HR��d��kf�0�O��l��?i�'d)q�/d�27M�[���@U�]����)T&�Zt��؟��	!L�Ĵ��ԟ�	�"G &{B�#��5yR@`��"|���%�L�K#"�+g�ȭ®�����W�)�܊�G #(��d�H�'0��(��G�&��0�<w�D��Q���N���
��	�\���O��fL+{�n�����U�ص�
@���I����	F�	�'>�
`K;	�I�7�N%�@��
7D� ��o�?S)��i!b mx��;�F�Z��
e�"�DTߦ�Y��,�Mk��?��
2��$	��D�`�83��١pF0aZHA���?9��&����޹6�`D��"4��	h���?	�;[Ѥ�X�F�b��� �a1 j��>Q�� m�,����_�~:���0��<M�1�[(iJ�P���P���*8:�8�$\��+9:��ɢ�M�ֲi����䣟^���bP�Hpv%
iz����$�O�V�hMy��$\��@�w��Cs�$��	��M���ip�	�Q�q05Ð�䝛� �[�z�^�[[���'q���D��9 ��'O2�i������c�j-��E�n�H�Eʂ�M<�9�	��\4׍̈́x��)�|��'=���	�c%���{�R�"I__�
�:�D�f����̉>�(����YKʨ8���I}މ��$-�)���M�n�]��ǜ�?��-V��'5��G��O����@Z�h4|��8S��T2��K�x��e}"o�F�D��ȋ�eS��B�I��'7�\㦡'�Лeߟ�6�ӷS�N؂w.��Z���F�U0N�<���~�.�RQ���4���\�������O�7m��d��6�S�d!���4M��I[>�١hJ�Z�aJV��|�恡�eM*��ْ�/
���KV69Sv�@ud��B`h��o5�`�3�
�f$�֝����[7�U�.̥O���%"S��
� M� pHnP0e��\#2���!�M�$�i�_���ش��^'I�2�O�4��i���|L왆ȓ{�>e rI���)� <kN1�wJp�(�O�}b�O��'��I&H�� �  ��   f  N  �     �+  ]7  �B  FL  1V  %b  Bj  �p  �v  *}  k�  ��  �  7�  ~�  ��  �  E�  ��  ˻  �  P�  ��  ��  X�  q�  H�  ��  ��  6   ` � �" �(  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3�����M[��хJ��x��#��+�$a��)i�<)T.�o��QՌ\�@��wga�<���4x�����KyK��jBD�^�<1�T���㕧]�_�D�R�(���D{��)R4i��	�`��>wܰ=D��#/$�B�	?~Dr<��E�T���W�T4@��4y�\Fz��HR�K�  *��[�_H(�"�J)�y�X���!�WDٚh�"K��y����<��mC�"f�d��C3�HOУ=�O�z�y�-ˁy��ey������ �'�ڄ����H�J���+� �.@)�4��>R��uG�s�~�{v"@�O:��ǭKS��H "O��*b�<��25cݾt�T�9��R��?�{����鳦
"�|�	u$C�_�D�s�/D�h!&Jo@����ꋻJu��o�n@a���s� �1E�Yp�r}�Ąʇ+=rI%"Oz�3`��U?���P4!�p��OL��DM�y�MX� �9�H%
08W�}R���@G�KbF �2�W�'�&Ö.D�Dò��RX����F@��\t��!8��hO�%g���X��}�a�Æl�nC�ɸ9�K&����Q;!&ՒyDc�اO�ME�ĥ�D)�d��.�"_k�ْ�mV��y�(��ȹ�E�V��%�DzrH-�MS��O�A�r�lڧ��I)��w�$,��"�	D\фɟ-<Q��c�'+d��v��gG�0���8-�� �(Л�8O>O�A�Ϙ'H`so.%�(��2�J5/r��O��&���}�Tm�Ot!�@HA2%N�k�%�>c����"��(x2C�	�f�.HH�kB�.�2E#B�3B,B�I�q�����	\L^�s����C�I%�e�g���Q� Q���yb#=�}r���q.Y3Pj-��΁�y
� �����;BL�Jp��|��L�c"ORm2iQ-���	֮�9�~E���TEy��d�OH��fiP3)O\�C�GܲY�80 ��i����)lUL�Ŏ�Tf�)A(��dc�Α���~�A���Վ!��`G��|�Ħ�S(<۴Fx~���
�
�8� ���D[��|��$\O�;s�	�&�J�Z�OМB)z@���'бO�ݒ�C": �|h#�	�I*U[�"O��b�A\�H6�mk�!�9I�H bR�x��)�� sb�]���B��k��?�b6,������ 	Oj-А
ܑ_��xar(&D�؊���#~���[��E^��6�$D�D���"�Ԉ��-=*�p�Yf(#D����˛,d怜�Wgֲ?B���3� D����AL1~p�h��4����/+D�����f��,~ucF-٪&
tB䉤=kʀ��_�ؤ��R�B�I*[!.@�.�#I��K�e�+٠B䉪!�nH01�̟]w����GL#O�n��D(7�D�T}��$�41�ȓ	�]�f�%h0�)���d3H���q�����fɯ�T��1����\��a�z�	d�M%:�H��%P=+��=��4>ay�들��L�'N�@Zh	��ƀ�yrD�VÆu��ت0�r̰W�ͷ�p<!��䍰�����Ar�KY�u^�	��M�O��a6[���h��@AՌ�����ȓm7FI�5 �?���c��Z���I�9��I[�j�1�c�#X_`�P�D�>�C䉟z�,,��ˀ�G4��U�)!{z�O<0��'��ı<qI>!�N�_ÈQ����S^�����t���'�6�KG�TT*D3/��ц	xY��؟�'��>�� Q�\��q�D�l��9F��#<ش����O�hiE��(b��[t!�� �
�O�Q�R��v�	���#����g�>��4��$4��L~���5��tu���`�9�N�'�yraݛ_�$a��Õ�UqB���I�����?i7e+�
��ĩ>�6�B+;j�+�M��=�P�h��Q�<Y�[7v�RA�U�&qð� S��Ny"�'�������;%�p[T��	j����'%x!�GJ@*Xmh��[
�����'�b��Ƌ��
fFMQ�I�SVV��O<�����F!+�l1��a�:�t�U*��P�b����
ۓ%���Ԫ�?��
�IB�L�xO<��D��P��� b��؂v�}+�)rf��O�C�I�1�rUPEԕ<����'��'�B䉥=>��тQ:�r����KN�lB�I���S�#R/.j��è_5j
�C��&	�^�B&Y7�D0 �#� ]�C�ɃJ`�gJ��)J�k�:6&�C�	"6�0lOA9y_��ئ-B��xC�ɫ&�j,{5IX�:F>|�%M�0�C�	�a��M��|�� @	͓O"��hOQ>��	!o�f<yF�7Q�� �Z����8ړ	�������Wu�X�$�pȄȓ$fE�t隦hb�ʀ��0�T��ȓ
nR�APs�&�R1��"_% i�ȓ0��ƅP�,FΨ8�$T���'����'�2��+�Iʚ1y��=�VI��'R\Lfa�	#RL�U�_��t��"E9�S��?�r��4�X���^.]��LP��S�<�V#�7tVE��G�/1�C�v�<y�ʇ:%Y�H&��ƪ�oVq8��'�\4o@}6�0��U3-_�A� 8D�� ����$�f �ma��m@a�u"O���dW� `vBQ�D!Jԭw�<�A�	S%��Y��	i�ʥ��Ky؞0�=��kIE7����F"�~\h�'�v�<����na �`B��.��$ f��M}Bb-�O~Y��͍DWP(�T)
c��D[v�'��6�zlЉh�$�B�9Ъ�DyR�'Ԕ��cIH^v|��ҏ:y:<X���;�������� ��[F��~>M�ȓt$�IP�X�&�� ����ze���I9�?y�}��)�&;	�	aYNj�h���#*B�ɕ\4���t�S{��iRg횄wV O�����)C�kT���!�����lѶ ��*O�9�� yp�,�7&S-<91�'��C���=�Af��2-���0��D$�''�tx�TB��D�V��A�(��l�'h.�[\�ɻ�&��o�ƥ�ϓ�O�Q�A���S��a��g� � �d"O���I M�R�	�FͧS�&4z$"OrD�SK�LP��Ks�Q9,�F�P��'G���D�����$ԲKN��cb�#d�HC䉦�\] rfμ6����*4F�<�,O�#}2Vo��h������%=:ux��P�<��Eϣ#4J��DZ�UF(���<)����Q�:�j�ʗ'$�2m;��2_�C�ɚI�$�x' �d(Qc�]'g��C�I�c��,[EÕq��HA捛�`NB䉜
q5�ӋY���Ë���C䉣"Q��;�.�97�4��OI��b����'�a�Tn�:��mu-.C9����
��y�ܚSTlM��-��+��Ĺe� 	�O����p2�-;��O�Q+�5������!�DG+S�*\0�EP0_�p餀�9S!��ڼ�8U�T��*c���0f���!��ȉ8�r���l�"N�����$�!��jf.	��

�7?X������!�D�@�.� N�#b���.[�`!�D�X�z���� q0u�g�_ 7h!�'H7^L�
2'����,Oy9!���Q��m�>h�^�0�k)�!�D�<[��h�A	�Ẽ��k�?C�!��A6|D�%[�*�29�.Xá�� }�!��ػvvl��ē����,I�!���!u��(�b}S�AA.:;�C�IA���7Ec�I�" �h�C�Ɇ;���mW�h� `&-�$hC�d�:��Q��S�
l(�]�7`C�	;7�8ɑ��L)XK�(u�B䉟j��AG���Mt�5��ڮB�I����#���d�x�9��G#-j�B�	�	AF���j\��hH꧆�
�B�	�x�YYQA���{��KvR�B�Ɋ6��Mׇ�u�� ��"�2,B�ɝF����a�'њq�=�B�7,�&���/Q�%�����9(q�C�I�V~K�.Ń0x����OE+��C� ����k 
_�������)U.B�=	�b�H��)x�(���A�=�B�I+%��i����M�dt@�c�>j�C�I�%O&8��̗��>pR`'_�MYvC�I+66%Ӣ@�*6�x�($h���"C��1<=�@**/W$����w$B�	�__��Xw��:�����^�uB��89�`�pV��e朒���65��C�)� :�I�Ç:^X�hq@��6!�� �"O0�2�>Pp�@���^=���2"O�5��6#�}�2ĕ9]�i�%"O��SM�6��d+W㏴�9p�"OR`��N�iΡ��ʘ�S@�'�B�'S��'VB�'���'���'��T�4�ހ3�Ts�Ѳ\�,�*��'�2�'�'Sb�'��'���'�$Eg����x`� ¶�X��'y��'��'�"�'�"�'���'KdP���Inz� �`H�o>x����'���'��'���'=�'��'T�HR����D����2B�"����'���':��'"b�'��'��'{�9J�$L�^m8�[P�s�̐f�'MR�'���'F��'C�'���'6�ty�jKW�����돠l���G�'�b�'���'<r�'���'P��'���u�B&<4�$�F8qr����'Ib�'�R�'t��'2�'&�'��QE�F9T��SAʴ�ݩ@�'�B�'�B�'���'���'���''<u�.Մר��cAķvK`�Ba�'���'�2�'�B�'.��'���'�Ѡ����F�N׫%t!���'���'���'Jb�'���'r�'�\�9 �X%GϚq���ʷ6�Иe�'�"�'�r�'���'���'���'����L�|^��BLQ�	R��'>2�'��'���'��-l�8�D�O�-��Ϡn�5J��ٷU��M���ry��'��)�3?���'��)����<*�]�r$���J3}2�d�v��s����&dr��$�@�%:A��99rh�����ЃK��m�'��I��?���p�fƜ��$�8�oƗ<o�xp�D�O�ʓ�h�� K%�́�Xq���,5N��  ��}9��*���MϻV� "�	*Gf������	���j��?	�'�)�2�f!l�<!�'���&-���$�)�%C�<��']������hO��O����A�Rc��B�k*t��2Oʓ��.���&�J�y�4��Vb�'Bt��M�+r^u��r!�>���?!�'�ɦ`P���h�p ��H�MD�t����?�!��<���|�1��O����W�쑉T凔*0��I���J�r-O���?E��'�`��疍Gc�����Ԛe�f\C�'*67m���ɤ�M[��O�6�2�k�'k���!�ᜟWH�ș'���'@��+���� ̧G+���h�X�J��C���c��πu3��N>Q-O1�1Ol��V��
Ѩ���΀��TH@R����4"��{���?Q���O���C�1v���c�`�z��p�N�>9���?QO>�|bѤ�$$� �ҥJG�ci؃2��!��񦥓/O��7O��~��|�W�s �ˆb���E<u����ae5�OBoZ3R�I,�p�Wh�,`mP�K��[!i:�I4�Mۍ�>����?��5�usq ԏ �E��(�:��#R��MC�O�:��χ�R��/����:h��`��\�l�����D04�P?Od���؟ ����Ŋ30�ȐӫC�#��˓�?��i-rL�̟,�nZV�	3P��p�0*�B
�qZw�,��8'���	̟��v�8�nZi~Zw���,�J\�g{:d�v��4�2��G�Iuy��DŇ(�CW�ϭJ��U�u	A*GT�d)�4�`���?���	���
A@C�Qߢ�JS�[L�	���D�O���0��?��E���^�g�$U�#I�^�|M������*O���~�|B��/T��
ñr��D�Z�9B�'���'o�O����I��M{2!�3L*� �(NA��9j���2A�����?	�i�2X���I���d�OT!2�E�5�rh��˃3yt�r��O�$M�r�h7�e���	�jE���֟~�){6}��ңe TB�PYEfQ͓��$�O�$�O���O$�$�|���b� Kp��AG놌�`)L�nZ�I6��I៼�	�?A�����I�杧~/�Q�oR8$����1��G;^y�	U�Iܟ�S����ɖ '&(l�<��lG(������'�E�,Q�<����
Pp��R�W����2�KI4(�ba�C�ս �B�I�
])U����dc�-V�~��C�ۙ�j8QҀּD*ި�ElU:b-H�/�q�=��e�7j��r��ԇ:纘Q�ۦhrn����(�깈@Z	m���s� Ce"�Z������6*P>:��0X���*���  �X�a�:��I�SGd}����-k6�b-͍3��(A�c�
�r�z��A��
���jFx�����J�*�(� &e�9����3r���Y3N�h���a���F��a�'H��nqŬA�$PTI�g*�F���t��Ol���O8�B��Ň=�0�%+��V�x5�������	n�I����I�/gH��=��Ҳ3c�|铊�Xq�����1�I֟�'�
�*aY>�Iٟ��S�e�^0��E7D H�� �(��BJ<���?Iwm�������A&�V�3�4.�tyH ��?D�R�@��Bɟ��Iɟ��	�?��5vk�9X��.e�XA�N�Z�n]o�����I4g5��?�~rN�U��r0���@e mPq����䢟����	埈�	�?ŗ'�b�'Aډ;��ԈG X����u�|f/w�J��2,�OJ�O>�	&Rp�@k�D&�H���J� SHKܴ�?I���?qb�ڀ���O����O��I�{26�١J��w�2��R�I>��b� ��I+���@������ �d�ݪ���@�_���ԵiG�e^"{<�	�����p$�֘�=���Tk1N~*�����o5��%��������$�O�$�O,˓z��#EROL���a�
�8r,����O����O�O����O6pᤪ�?o� ����i�4�V
��t�1O��D�O��$�<y��ʫ���Ɋ�,�`!��Rh\�僱�M;���?������?��q���p�YN��)�/7�4�;f	�;_��`P�x�	����	Ey")է}��ğT��S�/c�A�#�>r��2͒
�M#��䓕?)������{BB����?�ԚTσ�ڼ7�O��ħ<��*�|���Ο����?� +�Wt�9�F)�4�N`kU�S��ē�?���E��`�bןvX�'�N"`����C(�D�7�i�剷;������I���IyZc�2���'�\�X��oS����8ݴ�?���kP������O�5J��8`�Y8����J�
}n�q*�@�I,�	�����Ly��'�r��P���S�Ĝ�?���ؒ��Lm&7�+w��"|���@�8�#B	�Q�E��BRt�9���i}r�'��M ���h�I֟����t��p��^܊��Gz�h�>�Ə���䓖?I���?��5��cJ(�rݚT�߾h���'�p�P�+:�4���D�O$˓5&�����P�� �Wi�/�l"�i �m�=q�rR��I��8��IyR�K�2c�U#5�$�$�:Kp���1
:��Ob�$�O���?��OZB�:������z��W��ڴ�?�H>y��?�(O�L�Vo��|zW���F) �P�N�%)���FTH}2�'#�'������O��B֛,.LdJPaB�d��kq��4O2��O�P�r+q�������	��kB��G�q�f`��4�?A����$�O���6.���|z�+�INl����9��8�W�C�a����'V�P��yQ���ħ�?	��3�ݔ5@4�`bW�x���k�ަ��'���'"i�7�'��Oq�\cxj��F��C�9�S�4�(�ش��W�`���l�����O��I�L~"��(Y����djؙ:ꔡ�qL�M��?!Q.Z��?	S?��I�?���M�ʀ)X����L
�_d�0@�Ǧ��AC��M����?	����%�x��56� 1Rp�@��!�l�I��۔�M˕F��?9��?����.��$�O.x�ċ�J8�L�E��c��z�������џ(���K��N<ͧ�?i���E�_wP��X�J*"�@
Sd���M����?A��b!���4\?��O���O��� ��Xg����(߭ Ɛ4�iCR�G}p剦���0��~A��kR�SP�E0��)]T
1��O4�P�]jj1O��Ļ<i�2@�ZRH�&MF[u�X;S��h���"��$�O\�d,��럈�I09���P�E������%윒�쒮U�b����byb�'+ \�cڟ�ܨ���!������>s38��U�i�b�'5�O����O �q���Dț�v�M�!���@�D�*����x"�'l����ƥDj��'�0ً�h�;�!����_I�;�pӘ�l�I��F	i��OD�����{I1V�Ӻ4
�pIŶi�bQ���I'�Rx�O���'��\c���"o�f���`�ɍp�|��K<����?駋��n���<�O��ydO�m�\T��M޺d{�y�O*�$-�|�D�O���O*��<��T��8',�C��$��osJMm�ޟ��'��`���DBД�\QI�iU<Fi��Ч��M;���?y��?1����(O����J�IH��j"� �"Ȟt��9�O�����)�ܟ�I�ȸ1zԲ�K]^�؅�̥�M��?���*͊����x�O��'��b&ǥ=��Acf�_^�qdi{Ӛ���O���^�Y�pm��yB�'���'ar|J�Z�&;KƆ^�H�8v(�G��V�'�ʵ�P3�4����O��(ֆ����>6��I�L��$�i�"��4]�R�|��'�B[� xq D �^���>� ���d+�T��I<y���?Y������O��$�I�V P��ܓ7h��H!5��(���O��Ot���O�˓zܱbG2�.S���Ls��=	p(���P�����@�	^y2�'��a֦FU��N;e!�xv%�.�JL�oK�qT6��?���?�*O�=�ჀI�S	?6~�jF�"O�.t� ��� �М��4�?A�����O��$�0^f�d8��B�[��	"`	�h�ځ !�Ms��?i���?	�朇b��6�'E��'���㖧4�� ����CIb�p�K�=�6�O���?����|:���4���gZ�Y�rD0Püy�Č
���#�M(O,C�&�ЦI�	@���?��O�;}=�`!��c��@��O�؛��'!"HQ��yґ|R��6
U��(搓 �*���Z)V��o��6��Od���O���X}�[���RYt�,A�l�Z�Y��ʊ2�M����<�����)����0@����$�q�-�C~��arȎ=�M���?	�nz�q�U���'���O��	u��/-��0sΝ�HTFU���dV�1O���O��Խ*�����A�����ߠA5~H#�iJ�#�z������O�ʓ�?�����(�B�9�l��c'ǈ	��7��Γ�?���?����?���?)D�}\��*HX�sL�XdF0� )�id�'���'��'���O(�D�7-ݼ5���އrƌ�Z�!S9C;��O����O�bӬ���|Ҁ�	�8�6�;� �y��D�87�&�㯍�M�B�P��i�r�'��'k2S�P�I)h���&��Q%��!�H�����!XV8К�4�?����?����?Y�w7θrƽi���'`D$J�T�p�Lꁈ�J0�x��e����O���<Y�2;J1�'�?��'��X;��.)��[�Z	:ƀ��ݴ�?q���?!��/����A�i�2�',2�O����U�UOp��ꅀ͝LȒ�ic�(��<I�d��Χ��$�|�	�L�uԘ.W�1�\& ���'��+L�$Vz6M�O ��O�������L�c�Be�&j>��Y$�C
d�h�'B(%k��'��i>q���kǎ�V�1� ;Zp�8B�i�	k�j����O�����X�'��I5v��][ ��?��S���T$�y�4_=��Γ�?.O��?%�	��@��0@�(5��4ץJ:*��x�4�?Y��?�"&�5j���hyB�'��$�%M��ⲡI�16���*^�/q���']�)q;��)����?���M���Q�502-a��Iz=j�c�i8��Ň �����Oʓ�?�1v�p���,o��<I ��%��!�']���'m�ڟ���ٟ��'�����M[8TQ@I����D�=z������O�˓�?���?	�/�7u�Ɇ�E8y@�#��ʘ��?����?�����9O�-x`+Z�|��a�0.����+�T��FI��'Q���ş\�I}\扱a���(�gɖJ,������́j�4�?��?������(UF�x�O�Zc���1�_�rP!�z�h.���]yR�'�2�'2^�C�'���O�ͻ�˧t�JM�Aà�z���i[��'7��tY�}��~��O���O8���5���	�C�B��',�')�"ɑ��I�<�O;�!t��3'��3���"�0qH�4��d�j�m�ʟ8�����S�����9��JO�(��eC�9J�K�i��'�*d��'���<�������>`�$DY<	ؠ�K�M���EM֛v�'
�'�$��>(O���g�@�[����茍'}�ԁ7�����" g���I^yR���O�$H�/�f�V�FCP�w�%�5� 榑���(�I�_:r��ܴ�?����?����?��6hd@�$@�y�u�f�H�k}�4�O��z71O��`�Ik2c�\q���a��9DV��W.@��5�ɰ66�	�O��?�+O����;�L\8P<x,3��_�q������i��`V��y�^���	ӟ���zy��=~)2�*�њS�0�
@NԪfo���M�>).O�D�<!���?y�u;�h@�[�+%�t�4AN8y��]�<����?����?����?��s�8Y6�iHĩL� 0 �(�gB�	Y� ��Ja�j���i��'��\�h�'/�t�s�0�s�bʤ^Kjx)E-�	,�B`3B�i,r�'���'G��'Y~̢��zӲ���OL�8�A��:�U�yd@�piM�'����'�2�'����Éd>���ӟ��
V��VT�t��T��@:�B���Mc���?����?��ą�T��F�'���'���\&p$��,۞~O�T�"�P� 6��Onʓ�?� �M�|����?�/��	��.��u��kU5E
���K"�M[��?��a� !���'B�'����O�R�� (^xӱ��0T�.d	w�@���?)p ]'�?����4���O�ؙ!@�Q�;=�-�B0dTꐑ�4\p�E�i��'o��OE�D�'?R�']R�JX�$��p� L�Wv:���e��T��?�i>c�$��.a{���H
����U�	j&	��4�?!��?�$.P&}����'�r�'����uG��j<����Uv��*��K=�M�K>�����<�O-b�'�"�Z1����S%9oVA��e!av���$�0.�&���	�&��X�1pm��,7��c��²_t��M/�������O\��2��Q<S�1��!$)) .>Ca��E�Q��?�-O��O��$�&vXЂ�݇d~,��E:3RΈQQ3O�˓�?���?I/Ox���Q�|��ՀWX��lW�0���pW�QT}��'��|��'���[��y�j �|d\U�F]�:�:��f&�+݊ꓠ?y��?�.Op����G�W��:�n'U>��$�8	� ���4�?aL>Y���?)�@��<)O��	g�PZ��PpBCS�ܳqmi���D�OL����sR����'��d�FD|�E'ڲn�r�C%.�� �\OF�d�O��c��O�O��8X�ke��<T�+Q���,6m�<i��<��̢~*���Ğ���Ѻ<�R��]�
��u� �bӸ�$�Ov�B �OƒO��xiBǢ(�hQ@UcԻU�Ѳi�e0��u��D�OJ����&���	;pƨ�s��o;z�#.-�(�:ٴ�H(̓��S�O��g�8��y3�ȅW&vE�@ꐱv�F6M�O����Opr�H쓬?y�'��ᤇ�<QR���7���}�&G���'JR�'��S\�6T�#"Њr~*�"É��*��7�O|y�ΐe��?�L>�1M\bܫ�휜P�2њ�a���T�'��a{�yr�'�B�'b�I/#z5��I��;��� ��K�2lIs�V-�ē�?������?���H
�(�c�@�%��@�h$J�����<9)O��D�O��Ĥ<�2/�-c�)ߕO[\,�V�/<W��`�:D��	��d�I\�I��`�	�QN牧-��i/��X�\h��:z��e��O����O���<��ۜ.�OaZL W�Ӹ(/2��DF�2~��{�'h����'��O���3�~�>��L���Y�ʍF�*y��Ju!��O\��<���13�O���O�`� ��b�F7L6{rϚ�)h�0J�x��'R�-�B|��"�3�_�o`.hkv� C3Vٲ�iq前C����4[�������S����W lڡRn�%%��6L�9���'B�M��y2�|��逘}|��P���� rE�6z��ǝ�>7��O^���O8��g�I۟����DR��
r��p8�J�Mʉ������$�bм�"���/<�p��,�!)�0�m���	ԟ�AsM����|bI���ƭ�f��r��ڝH�ht�`lӒ�LK|���?���n=��+E �0��X�/2�E�iG�M�3N
�O�3ʓ1�`��C�s �l ���,7��mZyyB�'b����	˟��'���C��DB�y�$,@5ީ`�L�>�"O.�d'��?9���%a�tI1W��8R�.J�}4������D�O���O����O^��,�O�7�Ictrl � j�������M+���?�����?���R(��U즭´$Z06t�`��`��;�K��>A��?Q��?Q�t�>y8��i:��']�-�Q�,W�� P�Y��P��.f�j���OB����"\M�,X4�$`ӽHV���(`VT�3�i��'c�'0<u��P>����P��F�m���J9��E�֣W�(�b\bN<���?1�+�;�Ġ�<�O(��y�H0�0��f��"m��l�4�?���6������?����?I���?���5J��m��\������B�F����ڟ�����.�6b�b?]	��N.,�-��N �[�Uc�jg�P\�de����������	�?M��������Ъ
N�fEHQ:��b����h���M��7����T�|"�'ᚁ{��͉u�܄�̘�m����3F`����O��DR.pu����i�O��ɫ?��iՉ�rRb	��A��@�y�"W T������O����#KN�Z��׶ZE�̀�@zp.��'�l�x�^�L�'�|bB�5lB����aD�HL��ap��(���\c�Q�E"�|~��'���'F��'�@چ ����H�$�p�ۅh�F7��O����O���h��y�K�5m��5΅�	�@�#�ߞ;�%���|��'a�'���'"���ӟNt����\�4�ė�~<[5�i~���0$�������
�m��7R�<e��^!T%��F�Ͷ��I����I������`�"��l�I@?Q
;�!!��G��4�N٦���p��ڟ��	�^���g..���;L��j�CG�?�l(Iw�W��ѻ�?q��?A��;�0�#��iL��'���O,�48V�N�&Q� bS�E�5�boӨ㟔����u��5f(4f���`޵"���{s����M����?ф���?A��?��r���?�1��ڢ_��H�C��uW��mZ�����v 	�A5�)��7$i�G�*PK`8�U̖�m%�6mH��R���O��D�O��i�Oؒ�<,�վ2�-�T��,w��+e�	<D_��%!�"<�|*�B��5
M s��)c`e� Zѻ��n����ß�)a����ē�?���~�L�:'����3l]�(
���wNף��'&xS�y��'=r�'� 㑕B�� �C��l�8 �Kq�b���$&q8t&���Iɟ0$�֘�G` k�lL�q���u�ܧf��"?����?����d�=�M�vG�
8��y�ʖ�Д���.D�I쟬�IJ�	쟨�	0!"� &��Ҵ�"CI�|!����5�	�x�IƟ|�'q��"��f>	Ŏ��K���P�G�c ��:�x��˓�?�(O����O��d��>���$��'�z26]�"F3eEޕ�wZ��Iǟ��I|y��H�N���'�?��'X�b`�	 ��Sbbؓb�ϐ��F�'���ԟ��I�hB��`�D�Ov��G�مAn��R���-]�|���i���'_�	�}=�h�����D�OP�I�u���yGgՎ{p��X7��.,x]�'���'�Bբ�y��|�۟��H��.$����&a�y���Yǹi(�� 3��hyݴ�?���?9�'Q��i�ɹG�O)�Z !EI�4X<��g~�
���O� �B8O�O.�>�s�ICF��M"�8#;0�,~��8e�����̟,�	�?�"�OvʓR���U-� 2NT}�E��~�q2�i%.�ӟ'��Q�����|�DIk󌋌K�Ҕ��"�pV�i@��'#�7:�����OR��^�
!1 �ݷnJ��Ӧ)G�!5�6�<��_�S�?-��������BC2���B�r6R�(ed̎2�hTP۴�?��hֈ�?���j��ܟ�$������+H�
�̒=�����4��ñR����@�I��(��Jy2I�2?�������z!^����'��8�Ç)�$�O����O��<��ʌR�� ��l-I��|��H��|b�x�Iӟ$�Iҟ��ɦo�U��R���
�p���s��}����4��d�O��Or�D�O��A��ù4x��Kʤ[�L����"@=��;�o\����O,�D�O��q��3���V���h妃��#P�EtZ7m�O��O��D�O�T�Q�V�6y�h�
�OC Ћ��v��6�'��Y��U�T!��'�?a��>y�9�aEj��q-;t��A�xR�'���!�Op��68��b�IŶL��e*�Ù;��0��>��	��Eh4�����}��yڬ�	@��G�6�2�f��y�*��3��QxRA��&A<�k7C4F�jmICJY�.T��RE��x�+ӝ"���H#Ò�2il)+�D:Z���
� @�K���4ϰbf!yà�#c�K�^�@�!0��%l�Qq��	;82�Ԋ��� �"�#m�� �¦̪E�
�H��I�_9$�2��u�4�1�Ԓy�T�vDN& _�\���O����O����ź��?q��D����S���O����d�SM?�4�Snx���GPH��|)���n��a��C�%�O0����PD�!����{�ƹ�p�O~��@�'�b�|"�'�^� G���w�TLjRϚ�8q�$�:D��0�, �Rx��LW�v���h�cT��HO�Sjy�)�H;�6P�`ˈ�8@��K<��H�;��D�Ob��O\�+���O��$z>��a������7�:4&� Yj\7�����ط4.
("���Kx��ɐ�ַ԰#q@�k*
 �K�",(ԨP�B�9#�U�5d�Xx�ظP��O����	qfvE�� �m"����#�O����O���#d�,��i�$��#���|����_Q��c���7[V���'g�7'&�̓)���ry� �JQ�7��<�(�F99��
�..&9���L/�a�T�JND��$�O��$�~�f��uaųJ�S��/��'Ӛ,�U	��w�����̖�(O@�h�)��D���)˿� �x�Ĥ��m�(Q<.�J��R�D]b� U�~p�75SH��!�1h�NC�	�\��g+�y���#�M���D�`��3k@�T�E������'e��E��牄%q<��4�?����iV�M�Z���O^����V�R1ӹ&O����޵�(h���O2c��g�'�d}If��W��9���T�9����%��R��"~�I97��p*�C@�$��O��K�(�P�<E��'c6|�!CÌeWu
ċ6|�����ʆ� ����%�	,�n�Exr�+�S����C�*aE�6���KG�3���'
�y2�0:��'#��'7�ם�杩Hx�Jd*�@�a
uHB�N�!��g��`$�ؽc����(�?#>� �'��FN)v�sGł��?���8^�(S��G8��3ړ���i���Zo"X����J ��~�(���d���2b�ŷji"	`�$��4�4ȘCi1D��iTK�(:�j���-��*�� �HO>q!�Mӧ�#*m��	s�2|ހ�`�%D7�?q���?A��4\ϧ�?ɚO�Bh�3�5J,\���\;mhhyz���@Nt:b��;[����'��1���l�T1�q�ٵ =�qS�E�ٻ�ē-F@�z��'��#��?	�!�72�L ��Ώ��T0��?)������O��rw�!E���}Db2$MpSxI�ȓH����.���y�g�� �4Lϓ6�	lyrU�&o.6��O��ĭ|�.�پu�w�%�x�S
A1+�H���?Y�M�Τ���\�3��A��"�>�O�B�d!K�iW�M�g
BGl$3��$�)e�B��GO6X��}wK?x�A�����Đ�'M�#��h��Y�6U/`̩����D�"O|�B�-��M_��@k�9Y۸A+��'0O�٘4�ٔT��͛�+A�f�6�#�4O8D�K���1���̗OT�a�E�'�"�'��͐��U|�n�k�)G�\�d b���H��Q��T>#<!㥑��@��-�:U�0Ae�2����G�X�S��?9W�X�~O�4+���*�����͉s�p���?Y�O����O2���-E9~���@�%�佐�>Ox��%�O��@
�Q�p�ÏG�bΪ���ቪ�HO��HF���ǃ�i;�L3����l-��	؟8��À�QP����͟���ǟH;^w���',�9�0"�/M�%P����o:Z]0�'�p�xqm�:kra{� \��@�C:D
�;��Z��~2nR'	�4!*�'$��7�E�Up��S�#Z�Ѕ:��'�\Pq�'q����,O���<I5�S��V��*�9'B�"���]�<�׼>C̛��C^TY���ք����'��$�1^{��m��H�ځ��dI69H����{�,���˟��	՟��c>����|��L��$�d	T>������Ưt^`t����&�2p���K$��<��E>8��Ȑ�m"oIVX`gNکRP�-@B� 3R���b�\��$���O&�ğ'�~���!�1Ac����d�O���?��ʟ>h���yE4�q��� ��X��"O�q��B�~Խp�F�
���5O��'Q�'�\#}:3@W� �@���F�E�!P�/�~�<q3�L A�j0�Dɜ*7�N��ɕ{�<� ̜�E�ZAr#�
7򙻅��p�<�I�v|���6l�?�<3wb�<��dحC���ktW� �����E�<� ��s4�P�y���#vk� Ծ���"Oj� b� o	��I*Ԙv�,�k�"O��diĪ4�ThSGA�o��=@W"OD�#"+��]J�����2�"O`򥏌����,A�BZF�t"Ox(�����p�P0G�<��"O� ��L�e�jAq'�H1sC*��"O�U�N��MV�A���o/���"O� Z�JՓ �\A�,^�mC$"O�i)q�/d[*��F��$�Lݹ"O� !�A�x�����&E�9e"OF�!�A�1�D�/��و�"O�A�gOr��HE,��%�v���"O�A'���9��խq�� �"O�|���̑M��+� {�
lr�"O�X'��@�ごs}����"O���
�q?��	c�#�Y"O|I;�GO�F�q�����"�m�"O�)�)Ӻ#�Dq�f�O�հ�"O޽����L�{ �3(w
�h�"O.�I��o��9H5!H�Q���k""Ovŉe,Y�WI��c�f'V��ɴ"O*�!���|�Ը��dR'q�AH'�'������&n%�!����2@`���!�ѱs�m�R�'z�, �'�NU����:P
qӱ'��_D}���ɋN
D���[*:�Er�c����$�j;&=���S-d=�%d�yKޭh��� ӦT=-H��)�y2@+v�Z��T��Y"A"C΍(��"׮DM�H��OlɓR���ΉP1)YSOP�8fȆijy��(U��3��'H ȱY�_ת��(��Ũ��ҡ\ې��q�[�:��(�ь�>�0<q��\�M�6�r��E�6�r�W����>���9#A�q��U4Y�"=!c��q3��2�eN:3�N���cfY�a&ۼ4�b���d�i��|��I�N�z��1L���O�홥去k"�ơEs����lٜ]R�au ��g�fi�F��F�����T��Hqa%�C��=)2C�J�'�.��a
��1���S!%�T!��'�D����N�8X��� ��2�J�89��Ы��"}���xnpl���{�� �C�M�3�L ���&-����'"x��y�#@�&2F�1�ȁw�ԁ3��A�t��k&k�1]C��ǰ<���e��)1��K�r���1�ғ�p?���FR�eiP!��b�r��H6f7�,M]vx���K���ҨR*m���`��(�
\�v�V�V#?Is�M%� D�S肖+����"�֦�"�D�0h�t�
q�J�m�h�'�!��V�	;:z�:d��9�4��h	gj4�Df�dZ�bw�_�;<�AQ�R� ��*�+|�ƫ4%�4�@n�py��>}B�K�@"�E���#�����a���ClϷw|�4BDj�?d�㟴sVG_�vh��h�G�\�cc�H#��t(�V���cm���S��}�'v�9*�"Mw/��%�M+S�N0ja/�����s��)��x ���5�k�$�v�����\��mb_�^���C�k.>�>���	.	:ƽӗ�Ε>tT��Q�W�0ᐤk,�Ӻ{�'ս�?�S�|'����f��P�v��K�>*Q��D��G�}"�.$hz�EC�R�,���`j�,δ�G��`��ik�Ofhr����yRGJ9R��\21\�0�$K-�XKsɋi���r�$f���g�֕��M�"���ůo��x%E�;�����$�:xLݸ�O��!ђ|u-��&�
f>|���i;t X��ހ���K%nW�͒��D��v�BI8Х���d�!)X2_q�k3&��C��J�GV3_���O�z��`��杄H9�p4**]�!���x�6-?NF��I�X�4���Q֜,��e[�$�Q��Q�4	:��>aP ]�N�FXq�@��t��h���U·��I:rŒj۠�b�n#O�1���C�l���͚M�v��g��B��m:��F`����*��y�Cˆؠ�i �JM?�7�PA�I6�=�<x�qa�jp̉�Q�R��<�\��ǝ; �Q�']�<y�ui�%*�̈�	A9Qw�IL�p�a�`O�QKҘIVʆ�Cm@�;v���O@%'}���-���7�J�ig	Fw�<���&~�,X�P��2@�"���1hB�A���d@�>�@'c�T�U=&\d�I����5�>H��W?Oz�D��4����?��u�.h���V-k2�#�MF8�L.�)Vep���&L� #>)ϒ�)��8�B0��i#�!���@XH
��ۣu*�Р0� v�>�:����@L�<'�+����G����U�hQ�6��u�F�<���)g��a�N���3���Ӱ._������!N�`w�P>kJh{fM��E�K�C����F���S!����48>���-+�Jiy�nӲ[űO�<(�@ �G����ԫ�\l�ݨ��ɭJ�=*�H�v���	�Xd���D����� $�C�r����Õ:n��Q�F?O�)#���N9L���:�ŉ���%VΠ<��7�4}��͌���A.� h��Wg��D����	��O<�0�b9,��!R�Э� ��>����	�bnt��Ȗ8@y��S�P�p�0��.P�1�a�ȡ���)�
��Be�^���eQ�p٢q�2��>p^�0��Oj���[�!��i���C.a�Q��k��`mL(�gP�aB����igJC]�3��=N�H��K�Ȝk��Y jY�Cþsz���J;��2�X��Е*ѷp�J�{S��.5E��r��&=�&q���Щm��PW̾��{0�ۏNʓ ��q,�uG�֬G�J��"��$H�Ã55P��!�̇�r�t�=O8QP�)B,F��*����-�$��5��mK��ؠ`	0y2��A4p��q'���P4;�P��LZ�M��$�)I�e@1�d��"p�*�艗j��R��Qs�	B�Z�b�}��T�'�s%�ԡ�Rߟ��샫N��%RbJT� J�%eL5qA.�� �J�<	d��1�FuP���.J>$QdFL�`�J�s�-��aX�t�v`����"'�!��Gn�$I�cx�J,p�" �X��-��i�OQ>�Ҳ�_�IL9ڵFY���X�,M{ld��`��y�DY��%����b�#<�,��'$� X�n�P���7uϤ5	E��Um�	�a0pQ�DJ���	M��?�"或b)�D��h�$i3ʅ!���iE�`�)��CZ�Vc��VlC�Q�e
@B����'k2Χ^m44i$l��nY,$��� �`��	ӓV��`H�R�k��A�t�<E��ʄRm,��f���J��K�a��㞤��=�&�hgIE�pk0a���f��y�q��p�ؕj�� `I#�I%\����%ƋH��j�a�S�s��M��E�S
"\jASaD��H�b�z3��y�n U��H�� F�w��zP��O,�$��1RД���@�OٞM���ʞ`b�"IL�,�ɤz,�
 ��P����H�"Y�L��'}t�3Ռ��w���Fކx�
��OGM��{�{c����ol��eȫ~�H��9���0��I�����1;���ʧ]d��n�"�&�X�b�$j<M)
ߓn�L���ل]䈢竘'g��k�g�$o�Rq
�eX�_>�xp��Q�S���	^^���ې4?�d��]�
̫ņhNpy����+@Q��Fe��}��̦OV�y��6;�����ɪd �]�&��,N*X�Dkp��HH�5/�zP�欒�4����9�|,i ���6d���!,E����� �Zh&��a�ς&`h�iA2E�+_BR�;������� 26`����k�91��$��lp!a�/�O�ep��ţ[Ԗ(�VN/a���!�'�Z=�Ae��/����PB�dr�{*�rD�!�MJ��� �	�,�507�6D�dJ���+�>�C��X�n��<��*E�D�Lp��T>}҃ƕ�j]z({��E�<a�gĄ�j�c�Z������ix�����	6�FM�cf��r�����Wo��T��<�!מ!�Xyx�͟E���gno�'�ĽH�(�::�}A@NCD�P|R��D1��8�3��.9��є�	T�$
�d򸉔OK+W�x�B`�W��Q;E.��ya~2⑳u����3N(5�h�%�ˏ�?Y�A�?zcĀpUK����j6�S�S��n�L,r%
�&@�|�	�U��!��&4C�)	A"U�F+$�� �K�l@7��и��T�@VI&�n.牂m�����@�tX.��")P#D2��$@.c�2)�� Z�G�E��>]�"tqJ�t%�I�p���ё#R7w ��BS�@�+">1�R��p9#
O�5�,ɲ�z�'h@���{�Ή��R-e˲-��'y�ä �>0�(г�S(�h�:��L����k�<�pL>�|:�wԌ�sn����ᒭ�y��A���g�ص�>nY
���g/�ԍ�=�O����MjV&��e�o�pI�a�|�'BpH�e�'���b]>�&%���S�D�I�r<�  	�_]ܭ�W�	z�Je�=�O.�z�I2n?��Ys�'�D�RAr�����Z+B�h�ETj��ށj�|J?!#�${޹����t%�����3�P�,���)%吖o���J�� )\p�EMPZ��y�˛�mj~�I!ȋGo:1�ҋ���:0�ҫP<��ۢT���O�ɕ~�:��fVE�\���%�6|��x�diC�M���B't�M�Ģؿ+�v���sch�&0���J��9�) �D�I~��F��0���&	�2��5�	����� �x�Fx3r,�Y��ip�ހ�@!�b��?����Fw��3?�e\/lo>��g�+?�tx��ͻ��<1��_5���t��Y}R�S�@�\e#�u�F0Rq ��OE:�
�P�P[�bU�PӧuO�H��wP�ٸ�Sb>��	P:J^�xH>��Aր%:�%?�)�4�!�Z[@2t�@�# F԰LI�&w�0 A��r����C)�U�"��i�8��gɫ��8�rjX�e��ذF��=p�O���"'��-{�h;�N)��'���@7-id���
�!w�:�"B��2���7H�)��1��y� Q <��݂g�/���s&#'�7��(���gۏ{�r0p�(!��>��2\Պ� �K��x��E3��`*�O��Hp��> ��@'s�N퉃�D3K��]�D�Z��B��~rb_|rfH�=?����EP���T���f<qb@��n��J��I% �������'"�L(h�W�DыG���~��Ġa&�
4Ѧ����V�RU��	�pV��2���76�-��sqCˑF��EXR�=.�f��W��k dO�e����fc&O� :�3u�1U����uA�+Y�ՙ��[��1��S�u�~����C�1&n\{���zT���[Y��	��ƕw���(G������z睑)�.�p��n7����W��I����c���16mb�-a@�8D���'H�7|����,�,cD���/��$ٰ,\�D(���T>k���'yA�@*O0y�h'�l�6-	�/ $N$�O�%�����h���8�����'�$%��V����CM�z��ŐS���5I�L�"�w��m �/��`��iX�,ߔj2.�s���&p|�y��9L@�!h�6O��!G�����D�k��CG�%W��Ua� �1O�u!���,[}Ԃ��Z>�p�4Ŏ"��B㉡yĤ�����vZ����9"�CD�/,�\-b#�5��?����=P�"�ݥhG��a�_s<�;τ�U�����S�V �w!�1p%�!Ł�8�n��$�BNa�d �{r��p�2(��	N�p�sC��d�,�X�낮$0���C�
4 �YEx��kHdXⵢ�%�`�I��'����3������+�ͨ�i�4��8bڹ���V���Z����2�H��7���
,F�k�抮kd�#���>>cx٩�jD�&��B�d4�K!"�3ѭ�X�|cdχ�xO�C�	�lJ��(�.�'Q��WeR�=�tqˢ,��o}m��9�&���'i��>Ѣ3�*����aT���r#�6(��*��'q��C5-G�B����B��(����(�ӥ��K�aΓB[z��K>!�(Kn�OlU9�F3IAx��.;)�PZ���:
��٨v�&��0@�M(6��'j,�ve�35��i��A�P�ȓa��5%n�Rıc��H�F�M�b��)$Mv{@�R%������Y-,�V�;�;q�d%j���yR���1���*����Ł�nϫ���F�|~��z�%��<)eM:I����_�zLq��cDwX����֪*-��3h�	)�����ėڀ��@�.�C≩6>���͏2+���{���]l�"=a��E#_��bO�W�'N��Ѳ��`�͓��B�{��t�ȓ8 �SAc\#Uv�X�k���IQ���oȣQ��S�O�\D�r��3XܝbreƩo��L*�"O,M���ΤXfQ��%�qΠ%�����J,J�a
˓�00"skǰ+���Q�1�~���#.��:�j��|�*�(�U�r�^��ȓE�8��4|n��h�L.=f u�ȓ$�.��`�B8:���'F߬`_�}�ȓe�`A���P��H�Cf{�؅ȓ|���#:��Wl�*��a�ȓ��h���K�b`*I�C�5:*�`�ȓ5�����]�r�U�B������ȓ>�6Հ�&ژ�RA�����ơ��U;4e�7L_:��J+�Τ��Ц���!Jky,I�[�O2a�ȓ��`��偟�4�OܠQ�M�ȓf� 5��\&qx�PS�ɦ.�1�ȓt�n-����+�dq� &QLP���ȓC"��z��_�Jf���1I�!�ȓj~귊�<	
tBQ�M<���@+���6��}<�XU��� "O mb�$	bRa�Y�$KX���"Ox�摤+R��a�	�5);(�;�"O�ј�j�\p�l�R���%(���"O:�[k�+@�� q ȁ1||:�d"O�ES���*h�L�b)��0"�H�<�B��#�(��(�?%lmYĢ�B�<�V��:v� ;���x+���"|�<a�@���8����`0lՋ��x�<��_1Q��b��a���A�j�<aA�ʄAY�	�R�ĵ
���&�h�<��b1ιB�04,��z a�<�vo/'��c�&\q����e�<�� �!"i�Lq�K#?m=I���_�<�E�B(9���
X�G� (� '_�<��0!���i��w"\�8gb�T�<��P��c�E ��|򒤆X�<� �i��F�P�$<8T@1}-�g"O���@̅9@��\cIB�=La��"O��{�k>(#@�"��8�09v"O2ei���"<K��� �#��"ObA)3�@#^b�X�u�,$A� "O��(r]�64&��bӡ�\�"O"�HUoӀ���o�FE��"O��A-�N8�IE�Z��r2"Oȡm���`����&�vd��"OR�{â\ hN6��r�*z�*Y�#"O�AQ�_-V�6��%��$��Hj�"O��
�&��J����D��u|,�!"Ob�j�#��� qA�"�����"O0=˕lN9Eg�����$B�X\��"O��w�T.F�l�a"�!��'"OF5��K!b�$D
"�	5����"O�{��W�Go@��1�OE� ��"OjP����
S�"��"X4/Bx9�"O�\ʇE] C������`(�Z$"O��j��O� �g�=$�*�"OHŪ�m�~�dɹ���(<�"O�(X� ΍_�yb �_eV��"Ol�Sv/ކL���u��g�����"Oj����T�X�*xY4ʂ�H����Q"O8i�3�J�
v�	E�M�v<���"O�\Q��^	t� ��F�-,u~QA�"O��1��J���|��
AW����"O`9+���<�0���ߒYڄ�7"O&D�V T�n����K�R�J�"O��rr�U�v^A�U�n�<�1g"O�iF��e�~}`ԬJ.~xL��"O�I�.��!lT�!��$[f�4�"O�i�eh�1E�T��ê»Yd�H�"OT�P����D�H�C�� G�<�R"O6ݡ�<MF��lɒCA��k�"OD�#�r~���k�;1��S"Ou����tX �v)\-,B����"O��A׉!a���HU�<Pu��"O��ad�b� �p苑~+q�w"O�%5*=R��1%
&-�4ɲ"O�i"��/8����D�+�l�k�"O�Ać��B���� շ�n �"O|9AT�U�	�D��I�Fm����"O��j��-ǚP&�#Yx�"O�)�� *W�����DG�N,q{d"O��VL���AYd㚥t=P��"O(�s�fI5J�֘!��Kt��'�Q� �g+�o`:l�ǮQ�n�Q d8D�0A�ȗ@V(#3"��2���"D��!Aɇ�^�X����S�<�
s*?D�X�fg�o:��T��Blz�֏2D��@�IMA\�0��,v����:D��@��]�5��� ��"*wxT���|�#ғ��'����(ԔNtPШ��k܎�C�'�D�Q�Z�	:�`���^�^���'�&130I��<���H�Gƃj�Te�
�'Z�e���5lŰ0��]��X
��hOVв�Q���z���&-�
��V�xb�)��9<\�C�Ɯ�\��`0h�&C��%e�h�tO2�d8 �K�+.TC䉷"4���0��#�&��=��d0�ɓLSb���S�`3��Q�agXB�I�Ef�8�Z�Cu���R/ C�I�jyb��!I�}��ö�P�Q�C�)� 6\�d��l5#wD�g�hL��"O�3ԥ��6�T��ń�#tm�L�"O�MP�NU�5yT���=Q\N!�V"O$�@�CRRA��a�0!��6"O0P��O$F�<A#�ДR����"O���
�D�>=��O�!@�T�"O|2t)�V� \�Q�ѱ"O���1��@Mp�&�ɄD�*A��"O����aK�w"9�S���9�h�R�"O@��mG6}׊M�A��Fg�8�"O���3![>��([�.��E�"ODq�d�ː7�n��Ԧ@��T��"O^�JTGؑ
Yf�@�hX��"Op%9SIK��3��Տ	Z�� "O���6lQq�fQ@��� 	���"O�P�S�HN���[�O h0s�"O��'���q="ͱ"�՗6�:�a"O4%3F��4G���J&� ܖ����<�S��y�Mɝ4��٫��/'��"&�];�y�ʕ�X|9����"%z��T@�:�y
�I�ި�GG�w����y"�AE)��K���I
P�sə��y2ȧ'!�e��( R���nK/�y"`��E,1a"�.]� z&aІ�y2f�1Z��BTh��RqHh�yBlP,
����EtS�pX���y2l�n���1E�.7����J���yb���O��x[�)��8˲���G��yr��`BJJX��q�舡	<�4�
�':�Q�P�d[\��G�ٹ{/��	�'�t<��L:<�lAi���l��+	�'��)����vi�A 2f2b@��'%Ȍ�F�P�@��h�3jh���'��h��C-}"⍛�i�?��kc"O,��aѣ!�^x"U�T�)��%�"O(����8k��+s%�[�p�pW"O������0 *x���N�F�P}��"O��	b
D5VѺ���S/���9�"O��q�K>F�`� R/\��hT�s�x��)�S$c�&���b����q�K�r�>C�I�	���A18fm�U�lC��?F��hE#S _@�u�H6cv�B�IQ[���b�Z�0}x!���Q��B�	=q�	r�2-\ Mb7/�yc�B��
�@Zr��#�&�Jć��L��C�I+/�,t��Ė�Y�b���օLV�C䉬 �0 ���`�
�K��v:�C�I:�Cc�^�+/���Q���; ~C�ɑQD������ zf�ȣDiDC�	��2���	22�RԣA�a<C�Ɋ9�,P�U*)�J��D/[�C�	�2y6iQ�D�0qHd��
C2��B��L�:@�����,ThT��'D��c`LD�mф�K@N�'=h� �'D�d3�W�o���i��8̒D�'D��V�'w��<�׌%u��P�.;D�H�C�:$�&X*cE�I<��óE9D����:h�9�b��H*�i6D�\�5�Z� 4��D�6q�0l��/D��a���:�`��k��M��b��/D��y�(߃Dȼ�Ȟ�FD���*D�(� �Ƕu��=Ƌ��z���`,)D����`jЄ�g C�|���cG&D���A�ptd��S���/֔���"D�� :5@!��JeV���ű \��S�"O8YU���9�`�$�d"O��*�b[<V4�y��9-�僄"O��{c�� O�$K���:���IS"OQ+�I8T�׆��=�©)�"O@�0��N�vh�ɳ�E2{��]q�"O��P�4B(�b��54�|�z"O|e�r�!v�EɅ�$�`�x�"O�0�5`�- ���@�+>�"O��ܙ]|�x��EZ;�N�
#"O�U#��nŜHB�ƈ?� �"O� r_��(|"®�a�����"O���&N{��Xb�E:T��L{b"O�hSs�R(vZLAVC�]�t�
�"O���%C�/�D�����2+Ǣ��e"Op�s�	!?���v�5w�"��3"Oz�CAH�uͼ�����<N��"Opiyt"�\��A�>r��"O����і0���V[=(E�"OZXs�e�э/U�:��U�<a����`0!$E�(;*t����Q�<��M���e�&�l�[/�L�<���[�KMH�T	ʉ��-��nCG�<�'D�/��U�
S�<1x���aGW�<yf��, ��H�" �T$�|�<�vk��6���ʐ�@�4SEP}�<�C��	��)ڷ�Q,
�3�u�<a�J8��
���*M����p�<a�mǡ��i�ĕ�``�I��ih<�G�H#�)��	����S�ȇ�y�.��2Y�E#�)�|�ى3!A4�yBC�H4
��U+s���"lس�ybь1���rCO�d���+�N��yr9Y��0 /MW��Ige8�y��R+d�;��UZ��O;�y� �����C]׸H�
�y��^w64aƈ�f[�����yR�¸KƠ�R��Y��JA�_�y� #.�	`�o�P��AHV�O�y�Q�|���j�Iގ��aZ��yb끼�hcq'W�R��졑LX6�y"`V�W�`lKU�+S)yvBHxV4D�ʵ�3(5& S�%�fP3"3D����Ȁ T��2Mt�<�x#O,D�di�+�2ː�qg�/xD�%D��:So�6��m	U�#�\y�`"D��k���<"
��Ǒv�VhrfC"D�̸��L#~� �^7z�),D�D���\
`�\�p�HݱJ�2���(D�tJ@%��*ޔ���[���%(D�X�5lE�vj֊� ��ٰ�C)D��
bc�5��0�X�J̡ç�!D�L� ��9`�h(��&��507�=D�8+ԂѶ4��ua"��jB�`�?D�+��Ĵ��UM����Э[5C�	_kZ� �/иk��:e�9>B�I�45����F�?�L-"'���@,>B��8)!>,����
��Iw]�p�\B�	�v� �xW�F��@�%�0NXFB�	Ac`:��+W7ldJ��:>�2B�I
[0Ɋ�"�1U�VX"�N�,~J4C�ɱb1B�Q�.ץ]�f<�G�`JB�ɬ&�P]%g��I�Txhw��)�ZC�	O�PJTC�9]5L��M�&cvC�)� Nz�I��r6�iA[�p`�0"Ov�ZS�ЇH����f!�;Nr*q�S"O\�s�Z.�$�憑37t���"O��"��\c�^����_2�AJ�"O���e��rL�3/:(��A"O�(�6@	�<���3!cC�z�H�B"OL4���Z+�&����B�%"�w"O��k�dJ�Z����A�'q"�)�"O*P� ��7L|u��I���"Oސ��E��?����ac��F�|�<I0���f��ܙ6�էm�z|+g ^n�<��:g��S�,[�&�9����h�<)�ꄼ^,MsF$��3N�z��I�<�塖CSB�J��&~,�����l�<�a��(
j����r������GO�<	��ʠ<�@�f��.��1��f�J�<�ӈH6)ZH!���5h��r�p�<�a�>�.�Q���1?�e��Wn�<	W�؋>�9��+�[�\�2wn�^�<i��/B|-2�͚i��=�3'e�<�`�Q�9A^�[�j�A�^,"q�l�<��T�	 H[gS�4ri�r�<����,�8��A(H�S3fL��Yj�<�3`ό2��V�*�Z!)�R$">C��69��qĭ�!z)���W	�
[�ZB�+)�JI��٤H�F�:�����*B�	)�H�K�&	f@���M"t/�C�I�r�FlC&0�6��MK'&�C䉵{�9 a�&tq�%�E
�"qk�C��#eѬ��`��n��	�u��@�ZC�		]d9�v�Ԗu<��Y��J�B�6-���i�e�(��툥 H<x�C�	n���*���Is�M(7  "�B�IZ}� ��T�p�p��2�~B�	+�^5�q!E�
>8y�d�ƨ.C��6_�r�jd�۔L&y��J
<�
C�)	�؈S��^7IAcf�H��B�I2E�l��Ңwm��G㒮	V�C��
p]�����#�BHҠ!��C䉚ja��aW�m ����nN�S\B�I�0�``�'��J�rɘ@Ό�L�<B�I,) �`�#Q�Na��o�]
B�	�Z�ՠ�F�o��Ҍ�0'��C�	�"g$ęi������C�Ɇ�\�z�3F�~�C�E�Q��C�I2��� \'&Ъ��s�O��"OȃCN�Q��%z��sx5��"OpUyQ����~80��'�lE�"O�UiW`͜,z[��8Xh�84"O.��O; ����R�f � 	�"O>-�2-�x��8f	ݬ_��+e"OdY%iQ�Oi�}X��D�@8��"O6ĊT$�+
�^�Y���5S��'"O4N֢>4r�1��OEH�H�"O>�0a@-X�T�2�O�;�ͨ�� D�d8uI:H"�9ip�	�Р��e?D�<�#m˸�Ȉ�$��)��5R��2D�$�4��9�L��Űf�2h��4D�ty5��0+���`�A�h� ���0D��Ձ�C��y���	F��zUF-D���]�/X�eL��a��0�Vm)D�����*O��qZCb��ocf��')D����m�@���Ue۳,fbi�#,D�X�����t�4�
6�ґ�Uʈ4iE!�� z�t��Z0�/���7"O�+�����ı���V��b"OĉqF�%�N`�5�jɮ��Q"OH�R �OJ�dR#$�:1ɬ��!"O�u�H$v�f%�։Ɍ+�u��"O�Y8T�E�;aꄢ�j�	Y�DL��"O���X`�æ$��ru�M�U"O���H�W�D)�-�(cIL��"O�52'ʲe~f�S�L��8"OTe9�nO|M��d�5Ϣ���"O�PcuHQ&����ׯ�D�ܴ��"O�8������e��3�"O���-W�2��t��C2,�0�!�"O�5h��=�0���h�H�1`"OJ�k#��'T��P��8/и��"O����`F�=x%�'�3���"O� ��!��.��E��?B��-H�"O�ذ3)]�{��y��cW�.i0���"O�p����ֈ���4<NJM�"O����Y�p��८C�h��|9�"O�L됏ѐ`�B���ũP�>i�F"O�b@U���9��P�T쬺F"O6� ����^��)����%a� =��"O���(yZ��8$�ē8�d@і"O�4�@@ɸA����d��I�t�C�"OF�J �=*���w�S]�J���"O���4D4�����<A��tp5"OzL�f�+����� �+��""O�\ˢ)̉Jk��'�L �*��"OTEQ���g�=��c\�]�dI��"O�\���Ȟcb���A�K �x\b�"O�|��ϊWg�	q� B���P�"OP��.ӭ
J
��g�& �za�!"OVY���*aY���r�h(:""O�k��ڂb�,-�3��l%J)��'�RPcp.)7bɔ�͇}0�C�'�A!��/V��=rg�_ JhМ��'������ 5J����VI���q�'
L�����?���JFӑ��r	�'���j��!y�z��������'jԨFb��lA���Ph}���'�����Vp�x��fϦũ
�'�tz�M$���a�ć=`���	�'>^����\�f˸�y�G��_⾡�	�'� ��
��EB(�Ia�?K����'�ʌ nޠ�02��ۮEŀs�'T�=�1J��fU���R��'<7^�x�'�P�0F��: ��Y�
�2��'|�S��\t�@YE�*{����'�lPS��zV�e;R)#��5�'�j\Ȃ��:4�ui�*���i�
�'��*U	�\�3�b���	�'ϊY���TW�����y:t��'�j�s6�Wm șR�@T����	�'�F���lĮa8آ�K-�Z$��':$�Z7��r�P�eшq�dJ�'vR���Ono���5�˲k� ��'��	��f)3���$΁�N^����'�~D�F�Y�Y���C�4mJ�'rZTa@F�;!�(1�Ĭ�%>$�:�'������̻"����I+�J�'1��%(�$��Qq��˃D�4iQ�'�Q�RY�P@�I �:��T@�'�8� b�`��d��Ҩ2J�4	��� ���&��fT����Ϫ1T*��ȓ͐yr�BF2~�3��D�	�D݇�X"C�d$J�2�2�˫nKX��9}$�C�7tY�|J��]+5��͇ȓsĆ��E����(���ͪl?����P��4�5Q�
���.e���ȓD�2�I��	�T�$���W�Xh��k�Th�e.��&�t��0J�͌m�ȓl�0j�ʊ42��փ��),�l��@]
�r 
	6�:��ˆ�}��9��)��X���D3 X��u�N�,��ȓ�F�:sh�Mi|u��F�z6(��LO6��ũ��0�=��B�֞���(-2!�g�RJ)��bFKù]��x��s�|L{�=Ub=2��7J��A��c��@R!J�躍`�>�
�������aǯx�.-���ϲ0G�5�ȓj�(����K�Q� 8�̠�ȓkQ!�ˏ��J�RE�A�p���ȓY�*�DL�	��8�W�j t}��S��	�F#��
3T���&ư#��ȓDj�	�\7'ʄ(2�V��jt�ȓwd&aX�O�vE��O7eϐ܄�g��tҡK7-]68�	S.SY�e��
����?k�1�5�	nRՄȓ<�(�s���!!C8u%��L?��ȓ�6����ʹ��Tvm��^����ȓ%$p�����2("ԑ��$[ �n��ȓ>u��"lD�I.Mb�j�i�ńȓI��E{�A��Y���QAҬK:��ȓ!$�I;�7�A����g�U�ȓ�(C@*�;w˰8)t��_8��_ 	�w턕Y�t�h�+�L���R��c�	pg�p��lǫT����ȓ`$`��)�t�2у��-scr�ȓV�F��Q-ԤӄA5��L�� ג))4@��?�����ۓ��1�ȓG�ƅsGJ���*��S�1��H�ȓQ<(d���ƿ���ɑ�4��B�I���y�-���[�B�9�C�	�Yx��jT��67����A$�:M��C�I��d*�l͡\�Ҍ
V�=J��C䉲n(�ۦ�^9���*���4N�C�+\Fv��VK�(}�z�ز�ǌ#�B䉕j�¡	%�2-D�)Bb��Qݡ�$5��5B!��Ct�m2��Q�7!�$�';I�d��.'R�p�$l�
 $!�ā�:(~�!QN�lƈ�H���!��1�(\���!\�n���7S	!��hx�����(]B��-�:5�!��l����&͆�kx��u-��y�!�dF�]�<���Ț�MFv6N�=C�6B�=#V`%%�$�9`#n-�B䉚e��`a���v��4*d����C��	���tBŕ@��JT-V�aj�C�	�p����2Cך��V#��C�I�7�|0��m��r6h8`�S�MP�B�I>TD���'�/�d ���XB䉺"�Z5�� W36~����X�k�4B䉷a�BXa��}���E�bg~�i��"D�� ��&�l�v�w*@K'"D��Kd�%>ְ@W��p0���2D�$C7�R<�bT�@C�x��qS+D�TѶ�4'�����r�L��G/D�� ��:3,L�l�~� c�1���0"O2 !�Nt��
A��.����"O@�#�]���I3�]�!�T��"O�쓀�͇GF\��
�(Q����'�ў"~B�b�'����耕R8Jl�`�K��y2�ݼDR�l!G�0H�tı`.��y҉����h��i@�G�v�`����y"�[� ���P2��7?6� ҄�y�$�od9���ߓ5j�ҕ�5�y2��r=x"GF(�|�Q�ޏ�yb�Э=e�m��ϝ���!�� �y�nL8�eʇ
���z�P��;�yF�2�1e�K����'���y$�; �XuˇOPzŠ��Ūʨ�y"��q.��K��Z0y�V	+�����y2��L!����cRyA^�j�/ȏ�y��R�j��i��d�l���2�yb��*]F K���5]����ǯ�0�y�Њ���*��=P<���`���ybI��m�~A���نM����k��yB+G�lc2ŉ��;����AK��yb�;۰���h-.oTMZVG��y�(;)qL䊅k��16��6�yR*i�H,XPfժX��k҈�!�yb�U>V$Ő�DZ2v~�J�lؼ�y� �W�MtEvd3�E0�y2	3�x���kM�m�J=��HY��yB��~Y����ldT�C֢�yҪ;"f�$[���-`�~�)���/�y�	�%e���R�����Cې�yRh�k��!ɄU`f�PM��PyR�˜1k��H�C'::�����S�<i��̝b�@�*�m[�4Xl�N�<QP,Xghe �\8cU��T%D�<�G
��m�0���K #��@�<�Ǘ0[qx����.l��ړ�R�<��/V.#�^}����$=��@�f�P�<�� �z>e�!���2�( �K�<Y ���d9ށqu ��8�a�E�<a�G��I��1�
�w8��I�.~�<�����s����*� %�R��w-�x�<�r �qK�Ht�
�7�8��"O�<�p&���2�:[ �	��E�<A�,�`~=�s��n�Dȁ��G�<�s��a���F��e]�C4�Tn�<QR�=��P���J4�"!�)^s�<�3�V�z�U@@�ލ*�\|+��o�<ɡ�G8q�<�	�H_�R�9s!I�f�<����k~x��K" �j�:AOG�<��J�<x�����t(8Ĩ���<�A�P�>A��2�J���"��6iOs�<Aҫ�_=ڱ��E-0�l�T$I�<�u�ذ	%�zC-B^p�2�d�N�<	Wḧ.r��NM�ifY���d�<����A��鴅L�?j�����a�<���;Cǔ���O�<�>]���\]�<A�,^*1�1�#۴Ԫ"�s�<���M�D1|�+Wj��R�D����k�<�3j]���i
Cd^,0��t*�'OQ�<�r�H7D���� ��7Ţ-T��g�<a��оeʞz�@
?�8��e�~�<90c�)O�>պ&!��>=֩!W�Wy�<�&e8<��Ղ��ǁ5Dn�pDRr�<9S��PJ�W�]�\�Ka _T�<� �<��Ӝ3�d@�Җ/Hؑ�"O��@e(D�%Hi��D��9pA"OT�u�R2(���u�ۀP"O"�0�@@�_���ѓ��,z��h;�"O�Ayq�X�`-�p��A�=���b"O��լ~p�y#��*z�*t
4"Oj���J���W�\��\�4"O<�
�F���0"�Q"O���G����v�#A��2��D"O�����?x(܂�-T.U5"��"O�� r�hZ<�%V�~�hP�"O�ݩ�ІbF�bF��P,ޑ�"O l(�N�T�P����BJ-i!�K9��M��.
F�Mˡ�' !�Dߓ����R"��"�
��_n�!��]24��}�͹p�:QA��AN!��[��9��˙�A���\>F!�D_�[�@Q��-{f�`r@��$[�!�$R[�~�)��NgML �-��!�H�3v�)�e��.WH��3U�Ⱦm�!�\ o�ش���]Q6���녌Ig!�䗘�x�@ڮx���au!�\�5�	�ʖ�K����q��;u^!�Ė72���B �߫f�f�(b��!�D/C,z|��M_��A�5g:a�!�dK�B��5�F
Dd|ve�t�Y%�!�ć3"�RQ���pj��c΀�}�!���^?Ze��'Rw$���j��J�!�dP>��}�B��k�L��A)�!򤐟|<��IQ���(P�dg�1 `!�d2�&p3�jpD8;A�@?H!��J�w�&u�"f��X���q4!�$�@=\M�p.	#OL\##��8/(!�DŁ7�Px�m�dY��#E��!�$�11ج)����)S�������:�!�$�>:��Y+��E�gA��SD�E�r�!�Dɑ#u��6��)\&M��k�!�D4~�́
���D��G��l1!�Ǔ&�85�6���UAH(���@!�$ZD;��)ʄ�B��d�*!��&jw2�q#�L�J���00.V�U�!���1 ��#�E	yp!X�̙�`8!��F11�<�*�g��l ������m7!�� �={<`K�
�#3�����\z!�D�5KF��A�A�etl
��kp!�D��O�t@�]���E��-2G!�d]5\hPy(1m��$P#'�.!��� =�0U"a	ۚ���"�Ӽ!�mH�%Ѐo����u���4!!�ԩ"�H�˒���CLP*!!�DM,j͖�at�N8:�6MXvi׏n!��W6���
:�00Ti� ��'�ў�>�j4fG$r"��W�@�A�2�;��<D� ��G\Z�����0G��Hq4n?D��Zp*��r�DUv�_�1�v�[֩;D���b'R�	�B��T�	, IY�AC:D��ʱK��}���ܥP��qq�6D�P@X��s�R�n���0�
-,�!��)`���c �~�������!�DP7��kU���DT,#!��@�p8r�H�:4�������!��ҬA�ؙ�ۼɴ�b�E�5<!�$Oh�l��w#�)E�x� ��T?o!�$I1e���e� :�R���1
Z!�� "$��aް�T�����z��@�Q"Or�A�DF{�p{�`I<� �%"O�����H����PS �:>�)a�"O6����.��tB�/�uFr�"O�`�'�ֆSê"D�Q�Y+�0��"Op�*t���+)����&�݈"O�l�ac]�T�$���Gɑ_r��Kv"O^-×*I�q�q01�1\�جc�"O�xH%�)|	�����-���S"O���6��&���	օ>�4��"Ob�����9�$M�w��(���	C"O�Q���\�� <RP'D��v�h�"O0��M�G��Ȳ��l��*�"O�y��$^�ifjy{B�EԘ��"O���`f_�-�p8��GS���G"O�!:�">k{����&ϝr�Fa�""O��J7p��q�c��o�����"OH#@&J-NHH���`@��"O4Hu�@p;�Кtb�C�N	R�"Ob��"C�J�"T��&Ӆ+-���"O�A�v��>D��P�/Q=/@��"O�a#C�Aq�5A�T�4T���"O$yk`R�_J9���$ZS���"O��t�̜.�����<C*Q `"O.C�N>%n �a�}ArIU"OR�R	�3���$NG�(3�:V"Od�Qc��$wѰ��a╺lF���D"OԔ�䤆_ȬxB�� ��0*O��@3�n����F�]��Ld�	�'�j�a�h_�>�3dD��Xհ�'��C���Q=N=r얣P�T�[�'�b	���@v�!�qfY�#N���' ���"D��|S��,+��x�'�(�`��O1jk⇕7ܒxS�'�e �퍊g�(A��͒z���
�'��1�PDS�u,���\<j����'�fI�V&�9L����T����R	�'|�I�R�X6������ux���'5�ٻ#I�*�4��d�hOx!�'�FTZq'S	 n�QT��.d�-�'���!�X�$	�:���C~qa�'�b�Y��Jn�Q��L�=څ�'D�t�"ߴb�\�ـ�EO�`�B�&D��Ӗ�]q����bE:p��,�C)D����A0:�aS�W�n��0�%�&D��c߶%��\��	�8\ʹ�Q�C9D��(����r��dd��_�(�aO7D��b������e�O���1&k!D���4��?U'|��i.cGr58"�?D�`�$��	�M�R�T�r�(�V�<D��˵K¶]"���� t(��d0D���rə!$Zݹe�]XT)%�,D�X��QbaNI�ҋ�a� t��%,D��
�$B>z�"�{�Mh�,���+D���w�
	$RPZc�0����<D��k$��zZtH���)`Ɏ��Ӌ:D����ES�6X��)t�Q0�@x1N8D���#�$HD0� F�SK[���K8D�X	�H m�j�&ζf�4�pUO6D� ��� úlh�"�#� M �6D��R�(��C������d�b�<a��ͭpy&Ƀ��,)�,�`"�[�<�7���z�x�iFO٧h̠h(���}�<����XJ��P���J��Ət�<� l�6���"1���`���R"Op����%���xC&X�9��0�"O~�x@G��Up��HR�A�8%s�"O����I{���ӓ�A�S�.��4"OY��$�	P�Θ3 �@!jfxxц"OX�bc�tɎq�#�V7k��җ"O(H���܀K �	s�'a���F"O��2f��4j���� G=�ʥ�D"Ovɚ�hR5w�^Q� Ǌt�<��"O�rdܹXD����'U��m�"O2lH�ȓ{M�������H��"O��@�E
�E�,��%Ҏ,�Ṳ"O�Ѥ!�>�r�j�#FP���["O�t!���>V1�ؗ�S��j؁"O�h[f��84�|<��V y� �;�"O|�b��̢""�h��?�����"O�UK��H;;mda�
�#�&�җ"O|p��1 ���$<-[S "Ot���^���C���kI�xP"O@,caa�.H���)�Ʊ�8!"O�i�3�_/^-�uj0	Ӱas!"OQ��m��M�d̀�����|���"O���&��)���Y7/��%T"O4�I��X�t�2a����*.Qf\P�"O�1'͜�K�q���*w6��@"O�miBN��.�}b�	; �m"""O�%(v��RҦ�*@Y����y�A�8��0���3���U�B��yR�ؖxj]H!/��)z�0�	���yK�F��(���k̘iE)ǎ�yr�>}w�p��ܓV'�`��X��y�Q,XB���F77��m�ꘀ�y"ȷ7���>+&ޜ��N��y�R�0{��rS�߭3���31l�yB�	�F5ZЪ�)X�WT�| R9�y2���������:��0����y�8,�b`X��;f1��h����y�g�|�܀1�Ō�`8J�I�͒��y�'�#<B
�_��A��-\��y��ՙU怼*T�]��Z`[��V1�y")>����w�ǂj7hPc��F�y҉�=����)�(0}�`�w���yR�T�M����ш��"�6�p���y���B���yT�Z�T�Ц&� �y��kTB����S&�T�J�j�*�y¯�6 _��r�^���yD
���y�ą�:�}�E~�\�d���&B�I1n*Ҡ���$�[#��2>H�C�	1]b�9T
��K�b��M�X��C�I#@B^��Q�� (欨V��6!�XB�	�he>sҨ�	A�P2"�X&.�:B��1{�y���͗Bs�����'��B�I�v$���KȪ>��(�j�"�FC�	�P[��J�t�RT�O�;"0C����(����%<n���Ѻ/9,C�	7o��� b��;5�h0	��T� �C��'^k��Qf�%C�@pj�ɓɰC��34E�A˥$�
�R7��,i��B�I&H�J䈇^�h���I�v]�C�If0����	�Wb$���KϘaBB䉀i�(�*$D�k�L��"�A6)�C��2r^�3G�	��R��!!\�T�B�I=X��D ȑP�t6@�JB�ɝU� �`�ٜ!
�Z���8,�>B�)� �-�R��c�ܪ�n�(+Hp"OZESF͛�O��ZeC�51��"O:(J�G˻?�$��Sh�,|`1@"Or��(C��°�'E�6���3�"O���u��0k��a�CJ��b"O����Ə
Tiz88@�
���"O�4x� �&�*T�`c3f��R@"O:�1G�_�&@�<9��5�%f���y"D\"z�T20*ԟ#N.�Zu (�y�ɉ�\f
�p���!�d��%̞�y��I �@�v�$�v�rVdY��yBD��$����8s�>U�\0�y�j��BLj��e�dW�����!�y"�I�؅ ҭA�b�b���H��y�Ʃ30<�zq.نX�@�u����y���"
�527�W���3%mD?�y���``Kb��H f�Ju+��yr����ư�a'Әu j@{�OƎ�ykx�]�W���Y�CG(X�C�I�h����E�ą�������zC��`��5x$�H�D98���FZ^C�I�5����g]<�y�	�%{$C�	�;��A�� �~��1��;O��B�I�W#t�@���L��&yG�B�(a9QO�-+b�pa#�4#
�B�	+s��QT���L�Ц�LBRC�	�qS@��q��:K��8� Q�Ps\B��/?�X��g�R2t��D
�A*.B�"LW�4�s�ºt�h��B��N�lC��5�(
��[�Xul� Gm�4szC�I*5��jb�LOJ4�ABŻ.BrC�I�$w��afA�0Y4�p�M�/�C�I&v�p�e�O�Jl� ��W�C��:s7Z� 7j�+G�rĒ���B�I�	��ҢL�1V򴙂�o��B�ct���jC�+�����?K��B�Ɇb�ʉB��;0B�����MM�VB�I=^A��HP�L;D)�pƌC�� bH�2�/~�T���_�ZsPC䉪%?&�gK�>p��ʖ�%�B�ɘC�ƕ
�.�.O`t0�TI�;+0.B�IL���a"iWE(4j\�z���"O��{�0L��5[Ý<Z����D"Od����N�OT�N�.���"�"O���M�����#¨j�j$"Of�{6�X�d�xub��}�\8;�"O�XЏ_�EIY2���m���"O�Ī'	B?!7�a@�)W�6E3�"O����@F�IR���r�a��"O��Z�Ns�X���n�{=�Y�"OB=�e��=+��16��?'�s�"O�|"�(�(���1"�${<���G"Od݉Ə0A���&�'2n���"O�S�o|�E���X�L��"OT X�D�2p�x*�<d��"O�,�g�WbPd�Vo*<�5"Ov��s�Ⱦq"��IѲ"O$<��'��	@�hpk�K���Д"O��0��!k�`5k@G�ޜ �"O�Z�ŒZj�hx!�P�a��uC�"O��
Ղ.����jUN���!"Oĝ���lҖ��U��>�zh+1"O���Je,�l��h@�W�29 c"O��X�C�q���!`�
+C�ا"O� HQ`a#�JvI����,� e"O6(���M�<� g�'u�<A�"O�L�0�ڪew���,� =ba"OXt����qv �z��*0N $�q"OJ%���Lm��A �ň0BD�Y��"O�ي�EY�hE�r��d9�e��"Oh��A�ې{�Z@(��/}\]["Oz����8|c`���c��ON��"O�Kr��y=����j��G"ORMPD�K�#���3"�Χ	H"h�@"OPT��	��y*rh�6�X7��8�u"O�]�pa��:�%��0y�%�"O>��4-�(K�`�ʩ^r�eT"O��x�� CjD���� {pt��"O�$L�%����+X���h�"O���@�Y�ZR�]8���s"OP�J��YY�X!���T�Z�!9�"O� �֡�^��Dc���#{-:�x�"O��ien�|��4���3-����"Om�b#�4�ZL�ʕ�w��"OB\p�#�"�+tF�d�屒"O(�*"m��v$��2#&L4q��ڦ"O�	�䘌,J:E%�[��R3"O���!�o5:L��E�~��;D���d�?rD���īC�b 8�&�.D����?��w��,?&*�BvG,D�4�c��3$�(I�.Ҹj��P6(D���0�6�;�!Rg�}C!D��� O�=@��4���̽ �Xy�gO4D�(!�X�O�``W�mh�i,D��z�&\�����v�̴J��;�>D���a�J,QHN9��$&��<0�;D���g��B�$Z1�Et`;T ,D�`8�D�!.{�qdʻJ,�I�<D�8�q-a:8 ���\�KX q#/D�p0��BO�-���ۤ�4)`�D8D��#goJ%;��Yk�,�-Yt��S�3D�����%~�D��vmU�w%5y8!��B�XZ�D!S����"JՊ!���*G��՘׀�0�E���$d!�
�
�cE��1��|�g�A�=!�$�o�ȠG!�Tϸ}�cK0i!��&mǪ�2q��w�,9��C߶!�BC���w��k0cҚdn!�_)��EIBf�,���z&#��D�!��6p�`���.Ә]X
ɻ�`T)n!�DD�6-��ٲ �%=�અ��k!�$���j��6f�)m%�5�c��h[!��R�`4Z�ՃSj����_iN!�_����`䌖]rH�k���:�!�d֯[Z�@�ENpΉ3CB_�ee!�d&ppR���@&QM�q���gT!�d��2Ot��'��2qg(頰�^;h�!���H�t���C<;�P1�F. �B�0g��
C�I��"�C@�btC�	C`�ɚ6P�f�$�R%��atnC�I�d����G��ƅ�(�B�ɊƆ�B���ǜp� �)7 B�I�Zۀ��d�G�r,*TEN;#j�C�	�G��Y��,S){@�H��:��C�I��4��E�>X��h�5'F&m`�C�	'O�!�S%N7G���q��5#��C�	)ov$�9Ĕ�Y����Pm�3O��C�a���H=:a~(b$W_6FC�)� ���f�F�HfpBF��N�+"O����d�;�M�����h��"O���(���FΔ�9R��q"OJ���D�	����/�Q;ث7"O��9s��	V:4ő��$H��V"Oԁ�Woźyഄ[�N��`�aF"O�L��9a������t�+ "O�h8�ā1��T�'ɤc�=[�"OvD�`\k'2���T���0��"OvH�w�Fb��*k?",c�"O�QY�A�Y H5Ʌ�.Ș�ڣ"Oz�zS�ǟ�2A�B�����"OΡ�#��uX.H��&)b��y�"O��p��e��t��oٱcA^���"ODCt�l+�Q{A,��8���c"O���0��3w��5L͢i���ZQ"O ��AE�S�8����W���{b"O ���HN3q�B�֪ګR�.���"OTy����4��g��'�  "O����t��Jf-V1` ��:�"OȘ:tlF�F	 I���)26"Or���K��I8r$�c)Q�Q���S�"OL�@��;"�\(�g���"O�-(b��"|<��u�G�`���"OB�	W�  `�&�
�Z�p"O����e��<qJ	Z�E��N�$1��"OjiK��Ѣp��y��t!�I)�"O���G�R�n�`� cL$��x�"O8�b@�5&,�P��∗3ƪ��C"O�����Cs\ c�P�{�j���"O4a�G�#4�L��E��q��Q"O<ԑ)��U:7���F��t7"O�e��@ϓ/��ȇ!�Mi�]i�"Od���
Y�P�Up�U#. T�p"O� U��l���5.G?FŌ��"O 	!��#^����2�Q/8Ad�p�"O�%Z�*�0�G��S>����"O�萦��uʲA�f$�U%�a�"OZ�3#�>��\j��)+|�@d"OE�a�߽P�z��EI5:nՈ�"O�UzՇ��a%��@G�Ǎt�0�%"O�(!�Hv��qQa圣t�LEb$"O��PP �2X�=3&�ײG�"� �"O�� t#�����ď0�.1�1"O��-�^�@�q楓'5n")""OV��ǁ/n�p���_$bTq�"O�]#ЬJ����[QK��:����"OL�� �B W��x��$5T
Ќ��"O�ia"� R-�u;���yN<��"O����4YN�=�N�YPp�"O��14e�5�L	Bt�]�;��X��"O
�0�Y"J����dZ)�*�@p"O�b�E�x[
��t@����{�"OT��L|�pMA􀑫p���5"O�!���B�pŶ�aD�C 4�Xq"O�)G�e��!iـy2 IK�6D�|���^@�<Q�f��Z,I�p�2D�r�`һ'&� 4	�l*جy�;D��Q� ��^V�z��5Y�Xz��+D�L['+�*)A.y+V��C��X�/(D��T� r|�I$�[r�hJУ%D�zc��:�P�X��)2I�T��$D���nӷ}�½��ϲC4d����#D�h��1Jy�l���KC~@�#��!D�� �[��z�ˡD2a�D`�""Od�RL�	Qt�i���ʊ�j!"O�Ȃd�T�MR�= �̛:��;�"O�Bw��!����ԟ���"O�9wɋ�4_DĚ��C�q�����"O� ��%ӶH�����x)Р"OLQ�nµ-��
$#����h�#"Oj��A+I ��T`�k�&��e��"ODMx�[bΌ��V� 0��9*U"Of]��Ζ'5��=�’�%��f"O��A�͘�$�<�9�Ǟ;b(@{2"OJIɳ@ݗ ���䥐�YDbi�'"O��Ʉ��qs� ⓰>7V�Z�"O������K�+�R�J���6DQ^�<	��˟8\��/Z�U�U(sFRV�<	���-Hx�6�%P��d�c-�Q�<9�[g�$@��ػZwMP�#L�<��hތn�ؠh���a�8\
�\q�<���;�&QCP���:�"*D�<���ӟ[K�H��J�#�d�;#�A�<�d�̟� 9�)K�2d�BgZb�<I%C�R� �,�ˉd?��ȓYx���tg�<(�\�I1jܔ^d�ąȓ>5���j]� D����j�l��-��Qs��$�ӏO���Q$�[�1.�цȓDw2�8��48�����nJ,a8:Q�ȓE�*%ȃ��,eZ�K���q[�T��]�V���F�a�XM9B E�Eg�Ԇ�b���V�?K|
yS��8�H�ȓFlK�A��`�	)C0i�ȓ�Ҭ����[_^(@�/��.�	�ȓ,P0qew�H��@�{)ph��yt(��#S��hXT��ȓ*��Yģ�1�&��� &��͆���[sM9Q��3vcߥ��D�ȓ2�Z�h����*��v�$/(�ą�I� 	�$n�u��B`�؅ȓ^4hP@oߩfGn�t�̛+�хȓYG��c�c�W1��5��lo�ԅ�_CXmb�k�_�� v�؉W�����NZ~�2D�-L�jԚ��;A�!����@�/W6T^�1��K<�XH��M q�B/���҃U�p��Շ�$����T(�Sj�2��1P<)�ȓ_~�ʄ��s��P"�n�8Q��$��ET>p+ڪYh5�43[p ��ȓD�Աӷla���ӶE�.Y�|��a��`�d܈~�����Ò�9���ȓs�0D���W� !�sh�	E��,�ȓF�\�k_�?�fi�2*A�%��B�I<A^j���Ǌt2� �܀k�xC�	��ID�՛4�*%t��(�C��P�p�삎!�`�I��)\
C�I�P&���HۦW^8�2�ф%��B�	$s|��""ڊ1mLd�����{k�B�ɴ}�b=h婖;#;B���.Z8�lB��$~���c��)��bb.�5J�<B�	�U�ተ���w��)2nJ�}�B�-�te��W�J�d ���&s�C�	W����a^�C�n�3�耕 z�B� W� )EiW�u�*S�
_ e��C�	!AQ"���`Z�3�B���*2��C�I�Mm|� �'����]�ŧ+m�C�I�xy^�i��ߧG����ă=QhC�)� �x׉K�T�����P�$�l!P"O|+`_D^��!E�e$UX@"O�0!RM���<0p���H�@-3�"O��/��Ca��V��(B��	��"O��ʁ�Q?z7$4��o�O����D"O�����|���N[�76�\J�"O��W[�F��9+׍Iw�H�"O�a�/�����m�t*�ƍ��y�lBA(�аeY�k�ّ"* �y�+L* �����`:2܈�i_=�y"�0gG������*�j�As��y�ĨcBz���"�������y�� j�����d��M8� X� ˦�y��4��T��A�/KhޅС��6�Py2���9�B�QG��X�xEa��X�<��(�z�*5���x���3+�U�<їNP�Z=�`
Gj�~��,�V�T�<����:=�A�E�'/$i{��KO�<ѵ��#��ӗF����K�e�f�<����8���d�l�Ĭc��k�<	嬇T�p� r*!��K��k�<bc�U �C�*]/u9�xs�f�<�p*�(I�\bs"`px�%`�e�<�Ġ�-ALUs� �^�A��]J�<�N(�-C�h�QX8��L�]�<Y��D	E*|�{��-��u�H�o�<9w�M�~�`hґj	_G��X�]l�<)�JR9f��p2O�5h��H�m�<1�K�t	�eD�h(L�b�<�0$P/(A#�m�79�:	\g�<���NlP��Rs��e���@`�<�2!�>@�����O�.B0��N`�<���X'}D��x&G�%?&l��$_[�<���<z
���V�F	
��b"��X�<���7P���� �r컠H[T�<9�'�m�`����'H�}a��Y�<�
H#AI|�Z�#Q#!�. F�<�!@A�E�@$P����;�|����Wy�<�c�ƌW��Ъ&�3!Np�r�{�<�n-��9Y�fwt�F�Nu�<�Ai `�ޅ�Rg�`�@�ΜF�<���W6����\�z�����Dg�<!��۾p`����&V��U��MJa�<��D��`lՃ�?1�&T���Y�<�ޮv��l�d�#�$1�t!j�<��+�x�~s�m�*�H$�g�<��a�X�u�,/Nd0`�a�<I��7k�i��٨N�x��^�<�Gw�dQ��A�4�JOp�<��䀼B���S�~�X�
��`�<A�Mz�D��Ơ\�j]�%oU_�<)U���(��"`���4΢TB$w�<	��T�@�X0 `��.�u�x�<�@�]}�̸�G�Q̂�TK�<9�O�_�ȱ�(�~,n�a�IJm�<B�R7�ƉA�k�4�X5Iqag�<����;���B���w�"�����I�<��e�(N��;@.( X%Į�]�<Y�,8� ZVÙ�N�����Ā`�<AP���
X���&��0�"ԫ�"�]�<!w��=~v,RB�I$�&�[�]�<y���e�t��ՠ�#Y� �)@�GR�<�3%ԢT��pѰi^!M�JUѲ-�b�<�3ʏ�������^^nHɰGb�<� �e9�ݴ+�F| �+�3 =@��s"O��P4M%L�H%�jh�"Փa"O)��f��@�e	�3M��Z�"O­�E���̬Md���&L�T"O�Y��dI�k n4󁈎��ř"O�a��
Q��lp0R��.G��a"O���O��W�fx*nƋ,�UIE"O�1ʧ%��L��"�L��>����t"O�U�Rj*@H
�JD�I�]���r"O��U�Ef*Б��ͅ^|bX��"O�t� !W1 �bs�Z$[n䈢"O�]� HL�1j��5ɀMU�MB"Ozũ��/~j��h�52NƉk�"O���ܦ#���p�f�PG��t�ȓ)��q�/��>̴�q�L�7:|��Tw��ƨ��{�@��U�F�-,��ȓC������K"$ޤ{��@QM&�ȓP@�Tb'A��WƠ�"$��O�D0���"Ը�Ǝ.nNz�:�J�B���(lt�Gmj �wF�U
Э�ȓ;����th��_䑫 l�:I|���L���RK<z4�ڄ���5����w��[�iU�{��dI'�	�7Ѐ��0UB�&�Z.�e���\��2���G�z񓣎��R����n��/0�ȓ(^L��aJ8/}(��爻Y��͆�bl��H�;_�,���B�dR1��]W,�Qq��!*W����Ԧ2���ȓ�p-��B�e�
�����ny��uk�qp��ʆ-?$19��)q���[�L"+�i��g�#,�"|�ȓ<W5�MЪ]=�es#K�!Fz�D�ȓ;�0d��eF")9K��P�hh��z;D `B_�+4�ٚ���@��̄ȓ#����WeNA�:�� lM)IG����	�<�yrn�(YM��Ɇ�"�R���GTh<�B���8����n�F����	�:t���K� Y����H$j�蹅ȓa�����Վ}�6$�do  Xx��ȓ1#������A�}�CUa�ȇ�]J:pQ�]y�� 
�#��ʒ��ȓT(����&M7^@Q�b�X�������v����	��j��x+w�^�<�4�,}8J �L(t�隀e�r�<Q�'^�<���P`�@�$YC���S�<�e�#[Α���.0Y|kSj�e�<���N�a� iT�P��p��Ne�<!qE�AȌ��D�22�pۢʞb�<�gD�4}Ό3��((��%�X�'�E�T�X'WQ����Q�H����.�yr\����t�R�B�Т��N�PxB�i�8xKU� c� d���3���3�'>�8!�f�(�@ ��-��T��/��d�(6p�@��M��b�R����a!���MAT����Ñ1��u	�7tMџ4D�$�R���c/J[��y��C��y"�7���#�m�%:���Ѱ&N"��'�a{�*�Ȉ��Q_r���/���hOq�p����!��pFAsa���
	�!��B=g=�p�C �Ct�)�٥N�!�$Ȳp��D�_08��a��cw!�DK�o��m�tEZ6S�L���>7�!�dΨB�<�+X
B���t!�D���"l�E.�'*��X�,
�{d!�� �y�tJ�J�8���(#E��@0��	k�O�a���u��Tk�>�B��O>��A��Eك�A
dr�8D�~�,�o0>WQ�"|R�'�呲AK�Bj�����N�r�'i����E /?�-:��@:�MP�'��i�jP!:d9������'7��� XB\���1R\��8�'[O���?�X����<4�``���"o��y�Cj�(8G�IF���d�$�&E�p���F�l�J�k�L<RA�O�����	f �X��:_�I(�@H!e41O 7�.�	���'?��&F��x�ycP�*E ��� �	F�����)^��%�EH-@f��C�I�S���Dl+_�\4��M6?��C�Nl�����ݪF�� DK�<�nI��'�K9~kr�C҇@;e!!�Ak�P�d(�S�'L�T5s3@�<u�����TRN1´�)��LS1@��~�9���W�k�&l���,���<��I�.{bX��o2Y�X�a(P}�!�Lx�|���b�6QԦ�-L���s�yh<ٵ�.^H�\ZA�\��|��*M�<9�!�1���#c���'H(F`���>ɏy��.(�
��cCQ� T1Ak���vB�Ɍ_�J�QoS�Q;r ��-U�t�V�I֦�Exr�C]RZ$�A�>�z��2��:���y�*�#(P�rT�=;LX +W��	?�V8�ȓJ�։Bʌs<��r ���T��	d��hO���c��z���^�Y�bބ|bB�ɍK�RԀ�s�)�G�1	�B�ɷI��x[�.��2����V%�2�C�I
4�؈�r#��y&�8z�ӻ?�0˓�0?�2F���T�W,�}��daѩ�iX��mZo}�灊G�ޅ�Sl]
e`�dr����yR͚>y�����(`'6��!�µ�HO��ڌ�ɉ�3v:\Rb,
�B?"�3���N��B�I4ZH\�G��<f
�ࢎƌ`6�DK�������G�9!�epu�	
R���@���y"��#!�DM�"g[!谇����y�
�s�⠣��Ⱥ 9v�F��>4���=E���> (� `��.&u[�Ν�G�ą�7aV�	ENU��$|rB*S>"'����Ȱ<)�'��D�� d�P (��s���;���,%�d;�O����E�r�r �!�*R�XC��'A�OZ��+$�
����Y�n9N��B"O&a�'d��浻u���Z@LA@d�g�Iay���'P�0 ���;,J��t��$��80�'a��oϏ��*1�S��J���'l����#q]��͌�R��¶�_u��B䉾q�ĵa��Q�̌ɥ\%d,���v�xI�D7.u<����*Md�l�#������J~&8�7D�<T��7)R�~ԱO��l��H?��-;��+e�(I5@mㄊʠG��'�|"ŉ�/��`!�Kϵ�ޙR������$>ړ�~⅝�����QERs<v�߶�O<�>1ݴ�M�C�I���-�6��x�rTB�bRZ�������:o�ܑ��˄�h'��Y'H
�wyfC㉙��Y-��Dbb��l��B��hC|<��D�w����
�S}�b�D{J|j&.X���C��?�V�0���V��hO�O��m��'�8,��%�$�BD{�'pF� �ԏwʦ���)ۓ٬��'�j<�a)��_��$Yē�Gv�R�'�"�
5kX�Jw�`9H\PAi���y���Uz��yS*ʄl?m2v�(�y�)(!��a��̇cI>�f�8۸'�ў��� b��j��*��
�x�X��úi��	I�)��q+�O(=�܉�R7>	 ����8�	y�$�/�(O�N�;�p��v�E�`^@8"!�o��O���$��i,r�E�ͺG֐���: ��i=��'���?�����D��\V��Z2���,RQ�%d�!.B�&
O����],$��v���5�U�D\�hm�h8���F+P�&�x��V���{� ��;��I���Ө����dFI���sEm�۪˓�hOQ>���NL�3f�A�N\�Z6�ܛ�,�v�2����!*x
��6�vx�G�aZ!�D�16�ΖR�&�nX-�X��'�ц�ɑӖy0��*�
l���9<HB�ɓ4���A#�
 s��E�N�.B�*��@8P�H�E���k�2�
B�I'[�"��]�B�e*BB�wP"B�I3L���!#x��� 0l\�VC�,mfEi!,�2��H@���K�HC�	g�@!oV�>����&�W�oOC�87���oN�b����"DT6L�C�K�b�@�	a�@<iA�R�TC�� Lt���&��&J��-Թ�C�	pVH�G��$T�0� �� OS�B�I�|�����́)7�HTȡB�}�C�I�>��(���<8���JF�Iz�"Ob��5(-�<4zqm��
�,��"O�ce�w�T�c'���kf���B"O�'�Y�G��s��ǺNTs�"O� ��Ǉ�
� pv/\�
 �s"Oz�j� حr~޴����H�����"On�eh�B�&��sf�&Gv*�CR"O����mݞ	S''��(}j��E"OP}{����>��RLY�Po�$#"O�i2���!�q��V�:;XlP�"O"�(uA8����f��	��_G�pF{ʟ(�8ce	3^�Bm���G�>:B)�`"OY@��T!A��i��6}��9!%"OА�FbrD�&O�q��٠��'o��`�d��G�p{��D'H�.� F��!�dU$��ۖҬcy0��gD�[��	{?	b�铭2��H�&Js�0Ҳ��]ÂC�I8<�^\Q�`�w"t�1�+M�&���<�˓MR���P�G +O���p�10!*��?�TQ8�*Y�lA��"�0���ȓV> Q 
-"\�z�d�-�5��&�
�hV��W�F=����l�܅�_a��H6���=�ȑ�dA=
 �'�ў�|�Q�WS�}ҳjP_����¥�m�<	ҁY)X�!�׫�6|�8��%�R�<�܄&���`�����$1���Ye�<�g�Jն]�`i�"���k�(�a�<qU�U��n�s5�ӡ8��-�"A�X�<Q�S�Hc�i�'�R�!��	l�<��n-}�J�b�ƍ���ę��]�<I%�X�5z�AÏ0 i�y"-\�<A�R��hQ�7�#RHf�X�<��#�3h��8��ٶ=E~I�C-D�8����-s�q[Ǖ3A�B�2��)D�ةdOW����w��!�85�"�<D��p��R�4�MF�.*V�:D��9�Q�h'"|��&8�(�`�6D�D#2����dtj"��>M�yB�9D�<RWc2,�2D���\1i����6D�����N1Z��7�کp��8C7D��R�ą>R&�rv+X�?��ce�4D�� T9���X�&��a%ӠGe�"O�{�ǶHxN�k���w>>D"O*�1Tm
�\(�1M??%:��4"O���❘{���@�Ⱦ:��c"Oh�ӢmH�>z�iS��JC"Oz=��:SY���HT%*� Y��"Ox#��
`�ib�K��Z��W"O*B�o�	�@I�Γ��a��"O(9�R&��h5k�Nk��sr"O4�S����`���QΎ�rXR0"O^�(��ֱ{.�pp�-7�N��V"O�q�g�؃F�(XC��@��ey�"O��#�ʊ?���G�I�8i�E�6"O |�S�܂_K��4N�4Z�X�"O��hF oRj .R�C�Mh�"O���EF^"��Pmދ63�B4"O����AN�aS�<*��%2"OL��BV���y��H���1�"O:Iy1�ͽ/̖u	�,�}�P��"Oz�ae�ȄtɄ�1��V���27"O�|��k��@$©��/��W'�+�"O�Ò�N���",ˢT����"O
<)Sn��&:�#���(�b�,ψO Q��K&)$�[F��|��E3OX�y�f�2m3�\
����ޤ8"O�L�� �2F,j�:���!�m�"O&�����z*�p'��6>�-)"Ot�J�i�<_����B̾]ԴT�"O�����E�6!0-H0!��.5i�"O����5]!(���J]q��3�"ON�`���	G/Fd�5N�;L� !�"O�l��D�)b����kI�	!�ؖ"O�<���f$ �	��� x�u�r"Oe�G���5r)�&qBv��"O��s�(�<5�k�U�zڶ,��"O֥jF+C8]
��t�8T��ሱ"O�����B1E�z��1ʊI�V�@"O��#N�+_v�����e�lB�"O�UDjI<�IC�,�#'��$"Oe$(ЂWJ��D�F6;�X��t"O�	k��	G�N5��?Kᒨ*�"O�d�Ac�7Wp3�(�#��� �"O��Ї�Inꁐ2l��S��8�S"O"��т�9c���F�P�U����"O�B�ŭBS��w��8X\��3�'YX��g; U"��m�K�P����ڌB_��"O�Q�E	jwB��@��~㨰5�	�Ң��T!�: �t��@��?=uI�HX7"O^�p��Q�&E��N�?A����տ �#E��5��������썢 7k+ ('����Z�S��B�I�JP>U�7�֔9�(m9VLͫJA��������)J�flV]�剸 4�Ëa��Y��CI7&������&׀+�n����dZ�%�����¼N�t���/$�s�Bŧ+�ļ��:����$@?�L�-��-�ʨ��4��N�����NA��2�:�y%CV����	�,4o�8YB�$P6�X��		�h�z�Ư<E���}fJ��%�ҫ=Ӹ}ieN� g8e�ȓm��R'��<(v�U�`gޡU]v��(��a���[>���
�r���X �ԘQ��$Cc���U/J���ɵ3�Z��n�k&��#�@B32J<ኳ�E� �ZE@%"O}H<�`�ʕr�6�; �'j� -�q�l�'�`a�E
�A����ϒ�V���bֵJ��4P��C�<Q��XTZ(yU΁�Uk���G ����e��V�L�	�}��C��[@�O E��0X��<2�<���ED�!��B9�j�Z7'W'E��]p�'.,�&���֭wqp�'Yd#}֧� *�u�;4�:�@�� �ls"O�L)�9�-Z�J�z[B��j��3���A��F��̄�i��2�.�.R"�S��|K��D�.r����0�	2
��IK�{���oڎY���􇆎'��l{�������$X�=1~(	��[��� f�B�I�-çA�\��Ff��$P��\ÎT.g {gB�j�O袤�E@�<�����(�;�1�-Or@.J~����G1G�a��̚%VK�<[���*����`
EĴeEO1v��ʓ-�|�'�
��.-&�`)�� BOl>���h����(���f;��$�bH0�"#[E�@5��Q
�B	���->��T��s8�l"!d�v�x�·ڰ<�v83!���g��}
7	+y�G}b�2h��)�Y�r��,e1����	��,S��	(�E��8�s�$f������S%�Ksn�����1���D�5&ML�R��֯^�Oa��0��ú�8s`�P�4��q�2��"�:����1��+#J\��h���I�*�jE t�JBC2(�I�eY���@S�p�O� E��O��N�4y�z�Q�f1$H��V���y�Y�G�wh^	"�	�do��x�'ٞ�CTN�6"�C��
"��i���D�a3RN���(O�2#LY�!��q��M�;G~\!pϞa�����I�u^�G����SVYTm:�����D�[@Z0�=Ib��/%'��0�ȣk_�up%E�$��Z�19�i׆(s A�)s��ȓ8��E��i�,�p�X�",8���ٓ+Z����bkW�*�Ȓ����|��)-�r�'���w9��x� T$ʆ��Q�R��{�,X�XK�;�9O��+qc.N�١���N=� �֭=0 �"D�pq��30��p�kY8[�Ā�"#�NY	�>A�!ӗE��ذ�e� :s��� U1Tľ82����ƃ��0���?
�����/4�4%�?:d-q5G̓4�9�bעU����S�V�<Y��Q�V jJ���>8 b%y͟T�λW��%�d�³0���A���xN�,��'1b�)_�-���#PkM�jv��B�#F���b������ͺk�hѥz}�L
��@m��nή��Sc\�;T�%A`.MuAd��Ċ1'ԙ� �ȍ�?YV
߉+�l42$΂��f�q�e�����+F!G�<(#�Ζ�����D��K��M�G��9Q�>D�e�^�2��O|M�w'�%;x ���L	�`�֧~w�L�S'R�B V5�S%
�<E)e�X![�Ȁ	4"5����K�� ��7y0a�F�J9�x��4�����҆��/ٞiA�b�:�d�i6d�}�djޥ�C��u�v(���	~��y�+D�4	v�Ҕ#n}�3%���x3TbHdL:ii�`��8^��ka��1A �֝KV���	��i��'?1 �m ��d�@T�,�b��T�����,R�I�ɔi���+���$*�ːEG�Y�� M?|��mX��L!�Ex4h
��G|� �Vf ,SP���Oچ�qу��OxxST����y��R�]��%�#b�4C[���U;g�`� ;������U-V�c!FO�\s���䜌U��۳h�as<���@\d�'r:�¥@ݖa��0� �9���)F'C/\�A�O:�<�+J�����͐�|��9��'I�$�4=���OC�~~��0��#Dhy��O�[�8ԩ�ۑM��>��C��Ƽ�6�Ѵm�$�i�D0w��԰dn}h<��ne���p�+�^g�QzHp���	Ϙr�Z]��ڤe�|a玝c�#=��̄8붐�0�P���Xp!�Nx���@�Q/ ��| ����@�s�(�.�2��(_@�<("!�U��܊�n�22a}�+Ãd1�h� ��6��
����3�af��h�*(��̗�vd�#��c��]����`�6"���4��4>7���G|x�5FA 0��H�,&"(vh�ɕF�BG��I�+*"<S���T��]>;&���IEY��1�L�y`C�I�\�Έ�G��FTn��Ã�^��u�U��y��X4><:d��*��]��7鉨''�E� a�>h*���o�':����$B��^D{S��%Mq�3Ť�<m4�͓g*�Q�l���ܩ�f�d�Uːhx�xh�Bײ6�(���ߗb��+4/}bEU�,���(О�R�J�F^UT��r̜q���ӿzPB�z0Ϟ�hK^*D�yb'�<�4U���X?V�����a�A~�i�l_���s%
��j�mK��T�4ٴ�Ʉ=ȱ8qD4qM�IZ�+�B����Jf��s�J�HV+؄��"�@�ckA'��5�d��ҍ�-�*��$j�U�g�X�Np����My���ޠ`�"��#��#6T�u�3��z�`�feI\|�\K��O4��9�Ȁ�B�I�0?!b�GhZr�a��>U�$�`-DP��_�~(�T)�!�!F��0s��/8���B
�����@-&�pc�ĸ�B��Ń �q !�Y�2|5�'�K2�ɱ�B�1�]0pC�x���W��~'�xh��	��Z2�A�'Hh���J�z����E8P�`y	�'%0q7#ԓc)dqC`Ö�k�4�э�q3F)	��61x���O�� �@G�Rħ� X���])�@\a��T5_��c�'���艫o��=�g��,l�֣P)7м!�ƈ�+I�)k�%̈́i7�BC�;�O	�d�&��x�V����f�|�L֐��݃��P�I�(@:B�J6�l��?����͖��| �&U�"���Zv%}R�ͪG�;��|���ݔG�p�02@��TFP��
�q��&	����D�*�� ���INb?���)P��%�Ő]A�|ѳ���#���'������]���Ϙ'bB�z�י5�����״&�\�2FD-Td�9SO�_rUC��,2bF�<)�ĬW��iz&���H��[ ���c��Z'd�4ɉ��#�]Pɜ�4��eRF	�c�\�V�É�X�B��")�����*]�Z� `F�T����,m
l�
��N�1�i��a�%ڸ'�0��@#�,U�baC@�X�O�4P
�%�XH:1˗(���.O�p[�i�/Y�LH�Ç:�|��t��7���G��hu�bB�)H���xK>B�>� C<+����c΁v��Q��M�
:̗'�Q��-K�n.�ϸ'CD,kt���� ��7DK;�Z���F�q��* \O�)� }�^ԊSF�3�� p�
C�=�
=��o�/;`�O9��O$��?	���T�|��"M�1t68#��.��6\q�e#
68��A�ȟ����ŵ;��lA��/�zCq"O�,򒪝nkJ�Т�Z#�x�_��9�Ki�"��6��~>1z�MY<o+$u	i���q��F<D�̐��=ݨ0�G�5�Z,@���HiX�pR��y�g̓m0�Y�Kҕ!UT4���-c`�8��(�y��=e����� �d��d�L��Z�[��p��͙G��	/�9��G�q��Y��DM `��B�o�h�C��_��<�ȓ|U�m8�%��6�V�T�-+؁�ȓ.g�	H��W�8���J0H�+��5�ȓ{�� �t�
�&p��,�_�2܅��N�E��y	�,9e��0�e͈@�d���}7�y+���X�ȁNU	҈d�<����S�8�|#kS+;&��6K,�!��ߚ =�$���C,00���QF��8��Ɋ!Q�=r���L�^`��gݮC��C�ɓiV�i���M8�t̒`�5kD�9������ݦdf�xI�)�Hl��	r����;4����<�E/L,W)|���$[p9�W�F)��A�h_]�r��<I���)�z��W$֊mXK�ȓ�S�!�DY�
��y��o�rld�CN��p��I�Df䴻ԇ�8S�%K�dʞL\>C�:$�t`)7᜙4lE2�� nLC�%n1�	�逎O��t{��ǿR;,C�	?5(�s���B�'�|��33D��
�`^����!��|�1D�3D�P�$ Da�9�4��>k��DC5E#D��nm��0�����9�Ĩ3<D�l�����WpP�aT'�&aB8D� �FG3S ����Q�t�JA@4D�L���N������eU�t�tIq 3D��1c�@�r)N�Paeж2�^���=D�,#�џϪ�Yw�S�|�P�jC�>D��q��!Q�<�QQ ��ExQx�A+D�@k��J�.ٰ�BȠH��Z�(D��Y7�f� �p�6�y�h%D�xP�aåS�vaҕdρ2�D1�"D��K�oǔzx||�6)oV���2b'D� �4%:Mm�X�4q(��2K"D�(��aR�_"U�)W�]%4�g�"D�(�w���0(��yw$�%5Ɣ���%D��0��]�$�cpOۗ4��l��<D�����:�� ���S�ʃ�'D� �$lU�h5�8��I��̂U�+D��3�'����0�({�����g)D��!��-!l�0��Z?���;D�(�1��0>��[6M�y���Ӓ�"D�� n�z��_. ��a)T;K�� �"O���� ?���krƇ��<�Q"O���,�7��r� @�DH(V"O�E	����p>܊�oL�l��Q+�"O�,8����'��
�!p�|��"O i� �w�m��.K*K��)�"O�Du�Еv�-jǈ��k�V���"OB|QbX"Gxh�#gL8�x}k�"O�t�T�/~�r4¶f�/Je�� "O�A���Lz8����s�֬��"O ��g�ÐahL��ԍD?5��0�"O4aT_�E=���Ц��R1b�"O����(��0e��D��X��"O>�y���^�mC���Gü�B�"On��b���m��
�1-b5;�"O��i�m�MjX���\6��a"O�=��-\��q���p�NI�d"Onp����	;�,��r]6y�B��"Ot����'T<$�3�jO?�"p�p"Oz�k3�Z�2׾��4��'�ns�"O|��B���^)S�%m�9�"O��B��ZZ�)��U�(h���"O��*�)��u0T�uXN�P"O`��5H�=��u3"�?NJ��ʓ"O�9���
P�&4Y��E�;�Lh5"O�Z4&��oĸ=2_��E+͵R�!���� ճ���(���1��	@^!��
j��� �$\�H�6Y3Q�ܙ5!�$D$Vj�p��� G�*�3���;:!�$D�H*2
�K�Ys��
!�C�!H���sN�J��
V!���)]���a޳6��Ag�X�m�!�d�0=�!`���"�!�Ɣ'v�!�f�e�2!E�0�����K�h���ȓg�D��AF�Q��$�p�Z�X���yI.��!`´E1G)(@�l��2u�qj1��vU���Ub�(^ ����eg�x���D$��H *~E��2�N9ӌ �(@�0�V;o�M��?��[����$�jU��NF4��ȓq����f��Ļ�"��pB��ȓQ3^=3#�"Ymz�3��j┆ȓxL�-2������3�d��za�ȓC��q���HY�D�V�. `�ȓ,TPATJ�M��|c��Qv 0�ȓ3C(}��Cý\�VsG�Չ�"��ȓϮH�P�@�9UD� .ɆG; �ȓun����`�+5�H��%�%m�v���%l�rI�FΏ]��$��4CN�1�$�M��l����ѷ�ږOc
q8�B
W�hDzR�  ���s0-�g��;�-�T!��S���rgؼ�`�ȓj5P䠷�Ǭj�$�+ ��e-"�FCy�pВƌ���)�矼3���3�5qR���G�	��*D�����@�1o����F�9=j�"f����Yc�/-<~�1�qX��h�&.L5B��AN�T"��U.2�OrD�$nV�N6�����T����m�"cl`@$*Sh�:B≑vظ����*!W�0�-P?IS�<�d��pנٓ7
�+��O}���P��<�ֈ�"$,hZ,��'!�e��T�-��@�a(I\`@��B��Pe�"O�����S��?��
��m�0�Q��U�z%���~�<a1b�WD4��� 2�P�'�x?�bbY�K�����9��<���ީB:Vٚ��\	<� )���C8�@��Ȗ�_	��'ʓ����������ġX!�8��a>�9���R�VmxY1� </}��=��؎oK6��4�5�3� 
�Lي	�2���E#@����"O��J2fx4Ԁ���0b�m27�'��(s��9[�Q&rq�����Y��ZE��^v0���L�*�x%�ȓyHqS�͘-��S�͌�w9��$P�'҄�J�b��Y�,3���;��U�Q�A��1k��+D���h鬍��m^$F�d�B�� *���.�J���H
����, �2U����J�d?�TH��F�#��:s1��*E���a̵1�#`���!�	��(m�)<&��j��'�H� �`�j7J�O\��Ō�+Qd�H°l��el�)���3��$3!�ܮe�Z#}��0,�Ry#�㚪� 0�2o�Ny��Џh��;� ��`:a�TJ�	�4Qp ��Mt�1s� S�x�T�˒�G,�M0�|�'�
\*R�Z 91aKǣ/�h����d�]Pl�8�=���\�E��ҲJ��-�M�􉄛R��=s$��#+���"�Pd8� ����wI���F̡_�ΰ[r7-WT0WdA�~h�F}�h��!�Y��E��sG�vW~�Z���-,a�P�&�� ��O�5Rq�:��az.8zT�t�X�XO-���r��fܓRtrM���3����)P�aBb��ӥ�0-r���OZ1��	d�<_P��G_3L�)9s�S�<�� |�vu��g�DՄ &��N���7����7�H��	8e����I�������^F~�c�I �R~Ft���+��u�Ťv�e�������?ξ��-ª����?�d�ü�dEy��kX����V�k�n�YԄ̓�j`���:8�ni G�FJ� ��FV��X4M�9��↋{���ر`1�I=CHj���mt<� ح2T�L?a�!�� �(ms���zt�c�.D�Dr������<$� 舑��'k4�p�.B|�S�I ̤�S�����T?��'��b3 �O/��2%Lӳ~e:�IߓS�<)�&S�y�c�|:X�a!�܎VM�0�l^�v?��M��P��(lOI5�� Q��[g��,�Xr�����X@�U��y2�]$f���3�a	�@��߀h��B�lS�}+�<B�	'!�$��@'����5- 1�^ЫG��w��扙Y�(P3o��{��|�?�pm�d'�uӔ@���ٱ�"OdA���ߖ�(���Я|Y:̓���m��YiqH��Z��<��+|QV�0�Yֶ�#qh�[�P�h��a{B�����c������d��h�6�ۇ��l�m�f�xӘ$rE-�'z��8�	ߓ^��(�~dt;H��0��>AJ$
�bEb�$�>�Vj2S0i��O��a8�!A�{����! �/�!��W�9���!`2�^�Ǡ�%�r���Ɂ���'H�#}�'�F�Ca��i*�H�P�u���Bn�<��˘B�A8 �S;1���eGV��}	H�� �iz7�'�DLB������A�K@�/j0u2ߓT�@��ӧ�yRm�j# 8Y1cQ0��ŢH�נq�B 1�I %��O�kPM���O,	1��_��B�:V�X츑�I�5�Pr�O�,M;T�P���E�O�y��_4Lp�l��NXj!��#�J�e�$�Ol����+�� �c˜��d�(Ğ|r�ܩ�j����=�����hN<�J0�O�gG��b�i�m����%�dՇȓ,�HU�"��'pi`eJr�P(S��	�҈��G%tohmj�Q*T��9�R�i�(n���`�b�萅_�;�a���4z
B�Ɍ�>�@S=3$�9���8��@�J ����ß6Fr� ��8�*<�T�ɼU��+H��`�PJ?DD���dX�K��\��=BK��c ��L��g+!��B���2Z�����OlunX�BB9�O�M�T/
��"�c��ya!���|���|m
��߇H�����*W3|�g��B�����v<���%�I0}��O
�yB*��/G&���O��(G�Q������$?4f̘�dII�vz��j8��98�j�̻k� Y�� ή!�:��s$�;wtB�Ɠk�
�!��KAb�<��3z��Mb0��M�9D���1���^�� ��d+�,����T�1	��J��W:�H���	#c*$SŊO�u8�X��ҿ\�Q�"��&��4(7D��oL��2��*'R�p2�'��p�ǵŉ�� d�"��K��C'C��Q8�'W/�=�qB�9s:P��?��C�*=��q)�I� `��k,D�(���X�PmA%	'm0*5� 0}*�IZ0u�a)��q��јT��J?��
�h2�K��/��p�*Yf(<� eLR|U�%C"�t͜���h�`VR �Q:`һA�������Td#>�E�y���RR`%��=Q�-�]8��sH>� dJ�d	�>svB�^�a�L3��:$�Z����%q
��J��N5-a~r�� ���K#S�1cPa� B��&8dҐ�bE�(�j��q䓓pn�P��&ͫ.�3� T-{�)֙S.�
��U�Dat"O.mpA��Ҳ��B
�V~��S�E|�ȁm�/�$I������O�&@��`��<)��ݐs�Zy�#Y��>�8�	�\(<���%Yxx� E�� ���b�(�O�(a��'ǉQ3�q3 �-���d��Zv">��c�8i��s�A�:LN Hv�VJX�ly�B�;v��P��`�8��!.k��t�j��]b�EGĔ5�2���0?����4��W�Y�f���B��y�	�g��ۂK�:	Mx����8sB�y[���y���?�,����dt��ƩL>���//�*����Y�)�ӹ< ��UaN�1��)��l�������\�,I���0(*��&)?ʧm��d�P7TUʱB�<7�U��҆g^	M�<����$�>b>c� �vzSz�0F��)̴��˄�l�N���%F�`�pL���[h�H 򤄢n�@P����U�������6d�&b��Uy�k*�]�vH1���c&,X��	�3Q ���\���K�����&�9�|�Xqw�͍r8x͟8��"¶r���!M}�z�q�>;��;��D�����I tDh��kW�I�H�IF��(��	/_�2�CE��O屮�ᓪ Hpp�C�EĨ�����"L����a����'��#}�'%2��b�wcZ���[2g�b!���S���䛆oÄ��u�;���P��Ȳ�:,˖=��.�7���Y�-Yԩ��/ANl���O�.�d�؋��R�!�+~���R��`��0rToܤme>���ׁ],�ړ�1��p�����&�5YZd�̟�8��O�j��1��ʋ[�T35"O�8pRN\�{���D)�,y�AX������$_��Q(�Ga>�P��'�V3���(*R1���3D���c��jHF�	���Rr@,��>��	���,ƘϘ'aBx��\%T��X&@/����' �e�i��ݣ�ah[谈ׁ� �����'��1��Ŏ�oI|p�����{���'k�݉eH͞9l�9��"�R�$�'�t�i�Ʌ�<V(�� o�d?j4�	�'�^D�w�Ү�L���(YZQ��'	@�V�N#(��jRjY�'�V�񣝞n�I�W�O���B�'�B�n��q��)� L29���'s�y��G�.N�jע�	5P��
�'�Q��l.asW#U(]a�}�	�'mƱ;�ׁ[�������p 	�'�8�-�(j>�4+$k
�r��  �'��ł_B�R��Å�2>�0�
�'�L�)%��b�c���+��)
�'�\t( mō8��[d	\�6B&���'6���H�o�Ԕɐ-�xJDh�'���`T�2,�����3{MJ��
�'
��+0CK!}��W/[2���@
�'�*@
�H��������ڼx�~�J
�'O��;�k_,O�
��`���J���'kH��G��^��,���9`�Q�'ւ�R"�
�]#���4�ԌC��	�'��A�	�1@�(�H���SKଁ�''vܱ�]� o�5���YA�ܵ��'y�M���q�6i�Ӥ��H��C�'#���� S�8��	��.	�v�3�'G�A`�Eo�Ż���s���
�'�&QZ4��P�9�f��i1�)�	�'��p�GZ�k [֮V�^ ��3	�'f&)`+�X��ٲ�i��9֤4r	�'Ѽ���F�X�&��u,�>"���	�'[̔��c�Μr�
�ݘd0D�t��͋T�L!�p�ʡ	.9V�<D�����R�+�Л)R� cWm��y�@�����12F�< �LP�JH&�y�iH!i�x��S�YV�^�cf��)�y��ԛM��%H�6IY��y�"޶-m��[��4EDJ!��'�0�y���-�>T`Fɔ,Bl��	��y
� �X�Є�529뷢��Q�옂"OT�qUɵa���F��+����"O!Y� Ð��ia��G�y���V"OB���$��4�`ꄯ_-�Xa�"O\�K@��V� ɓ4k�5�%�Ύ�y�&��J�laa˔l�2��T��;�yB���w!�3bU�y�%�9�y#8��q�E�j)�,7F��yR	�ݲ@.��؈lY�
���y���| ��9�P���y�iQ�g��Deɱ��Q��N��y2h�]�N�S�E'>��}����y��T,=B:��WAٴY8�rL_��yB@����dj�&\:\s��w��
�y"�ׁJ�|t��a�9/+�m0Ђ��y2cъ-�~ݹd>xL0�		�y��d^�պ�/jHCFU��yR&��+XаQ�v���y¨�(),� [s��1cfL�y�۩�yb�)�(��vM��\!�y"b
<�|q�K$JҤ჋���y2o��mc�ɫ�� �r�L���B�y�$Q�[����OD(�N@�`���y���
�lH�5� �^�vlЁ�y�\ E�,�sA�E+� �B���yB�hP!�&���B��i
�y�aQ�-�����k���Jܸ�X�y��ͽ�hy:w��O�y�.ߺ�y2�/=d�u{U�ҲGЬq�d�>�y��\�|#P9aQ�֤v�j�H��ȝ�y�`H2��١��Hc�|��6��O49�5<�%9���dO��4Ok�W65F�U�,��p��8�O��9b��>`�f��H��}Z`�;i�p�uÀ�EH��)�З璸��/?Q6,�O?������1��01
`42W��-rј3��OQ?�㴊���d
u(ڨ	����O��=E���[�����	2[� P;5钬�hO��(��J��Q4a�6	�1�>Pj�i(1O0�S�O��%�s%��Xu<���P�H�H(O`��P'�<A�<�'(]-��b��ٲ�ـ�ĜL�\��O,4=�'r0aק���D�Jݲm�cL$HHE��AS�8��y��)&`�lH�I�< ���MĐ [!򄑮U��A+d��s6jtSacG�>!��%,u*)B&�: �u�����!�D �*�p\B�I�Bh*��q���Qx!�$A	W���2 �#KZ<i2�}f!����L1��O�L6]���zQa|��|�`�Z�(I����H��fM#�M��'�qO��N��O���l�TXi�D��m�����z�����'KV�Ж8Oh�E�T��̑0'ު(c�X���R�\"<�缟@�B.��ĉ����J����
)"M�D�����P`�32�x�����@��d�'�4+K|��C=�	�4C2�A��-ސs)n�c��L#W[L;4#Y�N��	1��ƻvh�4z���O��s�`��j�O�2h�"�<G|��8'�@Y����.!��{ԧ)���:�1o��Az`�aTD����,S�"�I$���Ve�i>�Ӻw� ��' �0_}>h���[�y"ۋ|��Ol�����cG� ]�Ze!�#�[L���
>wڍ{��#�: �"a��Z��d�s���-F!#�"O���	\�*�fJ��O� �"OJ�1��Å`�4��n(9�)��"O�!�Ǝ�=�Ļ�k�>j�ۖ"O���H�}��)c�JB�]Rě�"OE1�� M��R�c�#BTs�"O�%ۑ���a�e�#��`
���"OV��I�/r��aҦ!$
鲥�u"O�!�1�q|�4��Ǥbz`e "O� �t�e�['$�Q���+z��y�T"O�e9t�	c�1�D?Pnu�`"O��"�[�O���8ҁJ�QN��[�"O�@�(���ze��=eYJ�rb"O$�b�{���  [
TE�%�V"O�Q1��=�R���N�9j':h27"O���!��#� ��S-؁Պ7"O�m0�C��x`X�0vA�G��Kq"O.8��ۙo�����O�
�V�i�"O��2A�A�\���Š�5!�n�J�"O�ɻ&ɧ�"mHG 0�0�z�"Oe[�T�!�ؔ��ᖮ ���"O6�Kޖ��0)�!�!�R
�"O\�Qs ��S3��)Q��j�z,�"OhT���߮BX��jg��!���Ss"O�\b��Q������t�+����y�O�j���A��w=P`ᄥ	��yB��9�IC B�mp����W��y��Ǉl/(�)��mV*P�
�y��A�r�˔��s˒����2�y҆J�Z�θ#c*֪�䢖��y"�
�p��)E`��h��s�M�y�-,^��R1f^�����yR��=��#�`ë����'�(�y�G��1���b�-�5�'���y��_�'��8B���4 �X)0G����y�$��O�L�"��*A����f��
�y���`�LXjd�#�&�ҵa߱�y"i� Sg�d ��v�<�0%X��yr�_�qb�	1�(��lF�������y�̎&�hB��O�O�V��VH�0�yb�UK�~e�Z�B|)0�Ͷ�y��C���!C��A�< �p �DY �y��d ta��+�*l�U"��yrd׶#K�b��*rD����yre
F�XSl�4)��ma����y�a�:�5 ��r�\�hT4�y�뛪8�h��сF�
�Lܩ�H��yB܈Mr T"XQ;�@��F��yr�Yo{�a�t�ٙKy2��
�ydZO�x�+wY)8f�������y�-�/W4l{��T�=ؠ��7�y��h����n P��HP��N��y"��0�����'�AL��3���y�m�r��2	�j��SC%1�yrFV=nk�ac-X�l(�tAb T	�y��I�EE�P��iO"�Z�̄�yb�ӹEd��$��9fT����_��yrQ-B�j��1 �^��b0�û�y����F��s+�	M���j��� �y"8�,�3�@fp��8�yr�H0U��az�i?4����Fc]��y�;wL@��Ά2�$U�wM��y�I_%Z[���aǡ"��w!�-�yŘ�Z�A�g���!�*X�6m��yBӶ{��T�Bb�$.3�ћ��8�yBE\b<20���N�y�P�U
Ë�yb�L~(l]9B�1kH�K��Q��y¤�D�����Ñ{$��Jd���y"jQ>6��S ��<+jm;��\"�y"eC.00�����D�:N���qZ�y���)���X��K�C�H<���;�y�L�J�8��O2C�H5�w�P�y"�G !�Н�e
ˌ
ִH*��א�y
� ��꒯�2*�b0��ĩ0Q���"O�4z�!��q�\XR-Ύ6��{�"O�d���E���A�A͗�	(<X: "OP�Y`'΄E�
"F�~����$"O�5��ơ��jڊd���"O����B�%<�s�I="�Q"OrM�PQ���0�)�<��"O��a
֩�~�EJ�s���"O�!�\(q�T��GBa�	؀"O�e������ȽQ��{�aI��Pc�<a7@Xp( P���l�h��i�s�<Q�a0�fk	�*ٸyk��Ol�<��!+TX�A���K6\]ST�h�<y��38hl�LZ�F�>�Xu�c�<)���3B`����� ��1�%�x�<q�jܞl�Z�7
��b�ↁ�o�<I��E
P�E�t/߲��%�eBt�<1��,K����t#�X��0��Cy�<y%KW�>��9s��
g�5���Fs�<	����c#�I�%pa��Z�<�MDl
K{i���L'>�B䉟� h@`a·PIz�YcLG�/2B��I�PP�amb���Q0F���B䉲$ʼP4��!<Fڀ���5*�C�I8�|����*+$�����0?4�C�I(�<m�!C݆87`�8��_�!��C�	9v�2�� ��z��Ł����AϘC�	�"�X�uU�K)�1Y�Ƌ+zC�	�(Z(Uq�����)��aC��B䉮OV\-`�MM�#�X�`A;y#B��N�TSa��l6�@$ *V��C�	8 F�ʆa7aP�\�%@:F�`B�I>.41�l�?!�h�h�@�q_DB�I�@=2= a�\�7���G�TdTC�I,rE<P�#s����g�&�DC�	�i�ʑx�d��r������C�	.�88��(�7{9v�2B��*)�C��0A��c�ps��0&��2ޔC�I����6��[orQ	�I85d�C�I�+Q*ps��� �(�@����VC�	�	�NyEE3dS�iǡQ�0�VC�	p) ����8J���O*Z/8C�%�>Y��H1����2,͟p�C�	�g��Ԫ�Â&D_Yc$˒c?B�e�*�Z��F�e	&y��a�B�	�.=�`[��1B(D�����#��B��8S��ShҝR���aq� "��C�	�fx����,��{��m�0jCϨC�9�"����V�*�����(�f[�C�	�@�l�(0d�'.���e��I�|C��x:<�0�]�r��� b�Z<}-PC�I`��a&IH>+��3SgY�edC�ɚ�`�2��1T����J�hAB�:nl��T�,VӒQI`�V42��C�	��t0$L$�6)0�T
3�>C�	�#L�b�֭\�*�ٰ��yXPC�I�|�4;��(���A�όZB�U�2"��'�j�"��+|��B�I�U� xz�i��f����/��B䉣	�$-�Dh^ m �Y���fB䉺Q�hxp���R�̍�3$�17 bB䉦2cRA� F�baz�"A�P#�LB��'Re�� E�`�8�B��-~�@B�� ~b�M��'E�v�Z�HFoκ<�B�)� ~�*��IvH��Y���kK4ĺ4"O,�!���@��h���Sa�%��"O�]���3zh�(jrIB�"W���"Oƽ!#�.�,x҈�'V&��hB"O. نEΩU.𻃇�H���"OX��UM�yݢ�JV-�HI^�5"O\ԁf!��Ln�0*�0�v�R�"O�h�"�h��֢�2*� ��"O
E� 萫l�P�h��U]��h�"O��W%��k{"ɹR╄\�.�0"O̸# �3W�,� L�P����"O��@"�!gԭ[�I`v�i�"O��0f)�><:S��W�pb"ಶ"O�`��"��*���	V	��&`j)3S"O&4sw.W�'��0c��[P�"O�Hi����1b"��#M�L�q"O��B��2lJ��/D1hq�s"O&]+�����-)�̄4��P�"O�!sp�N Cb('���M��}r�"O-����$Q����
ϓr����"O����(�jEp�K��q�"OބbB,]jE�ř�$�=7�d�	�"O��#釖n0�IRV.&��h[1"OJ�����+=�h��c#���
�	a"O�88��R��i23�Q8h��V"O��w�H�"Ȉ*��'�(XU"O�*2 ��#�:�9d(S�Y�Us�"Oؙ�vcZ�}�VQ�W��3.���$"Of|���K���P!�90���"Oe��S�8���q�o�4%���!��!L9�!�V�V�S�.I�0��r�!��R9�x]����2��P]+ "O��Q��N4����ek��v+�8�E"OD��%��>�~�8U�	�wpē�"O"��"ω@x� ���_�q��"O\!��)J�3#Ș�	�е@2"O��7�"��s�Ć�S#؅"O�T��m�|^�Q@�L*3����"OPm�Ɣ1y9\EB�,G$
v��"O�hKsJ�*a ���LI�d�80"O:)ZC��`�>�alY��X(�"O�D�e�IA)���aO�=�81�"O�1�M��p�I��ry"({�"O�bF�S�g�.Xۄ�K�����"O y����2��t���]5!�t��p"O��w�l���G��[�U��"O�}��	 �0B���舼JVN��"OQPBl�4}�ب"g�._���kg"O���vޓ��eyC��?���9�"O�t�$N�)�$� �d !��Ţa"O�ٲ��*f3~M�4�Йc���K�"O��y HɠE�t�	��V�\�8�"ON��9t�Ash� C��y2�"Ot���$�`R�[C&߻q~�	�"Ol��ȍ�g�Uyp'̭d��x��"O�@�b��	�Va��'�6}��T�W"OХ:PCR�(��� GC1N���;�"O�[a
$,E���V!a9R��1"O~�z��@�O�Y9U�Z-�h� #"O�	����nn	�҃�<Q��<2"OH�@ 
  ��   E    �  �  ++  �6  ^B  'N  7X  �`  Jm  !x  i~  ��  �  ^�  ��  �  (�  j�  ��  �  6�  z�  ��  �  H�  ��  9�  G�  ��  3�  ] �
   � @# y* �0 �6 9  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�ou�!Dy�'�:� Ή�B�\O�|�����<a��$�+q��@rsI�E�f�W�]�1O���$���R�W����FޜO��'*(#=�O��)1�h�Z��K�`)����:o�.�<�J����<4���y`���`KR5��O��Dzr��`S��o[X�JC �+�lԛ�#D���5�^;Ki�e:	�L�� 3 �6D��@C�>y��HRc)ȓD�* �$?Oz��L�r�:M�\�H�| ���� d.���'�.���Ǒ����r�Hp*QGz�~RQ$X�E L��]O	�fe�y�<Y'�J�oW��`2m�V$��s��Any��'**��%�T�ncL�@���h���'���!#kB�踬�@ˊ	�2�#�O��G{��4F�R��F�|�Sm]�y2��6u��	��݆i����y��K�eb�#�-�b���q�����Otepa����+TJ y  �0��rL�C�I�t�@m��'[2H�U�LQ�!>Bʓܑ��|Zjͪ<\���,B�~�!�a�B�<��F��@��4�S�{hh����u}BX���ڴ��'4��'o��e�f��;i�(1b�蛞09����Z��� ��x	�aqP&�3^i^�Gz�D(O�e(P���0�2m����
ba���"O�mkF��f�-[����gX~��"O�Q��gX=L�(��kL�*mA���[ԟ�?E���P��,A��ޛg9(\���C�̄ȓy���C&�6��[�M:_�,T�ȓJ����X�%;4�҄�B�kTL���	|�$�8v��Y��l:n�뀣�;RV!�$ ֒��O]�6ě� �HT��\E{��� �QZ'���Ԍ����<	���"O,,�p"T]q������^`"OL�:���\�Pq��@Y)u��x�&"O�m�S�O)t�~T�%IM)n�-J�"O@|�㢇s���ʡ'K8IO�ܸS�'b�O�l
&C��~"��ᐙ;�fY���	4$E������}��p�'l���L���<}Bd!##,h@���W^`򣉒�yRN�C�y� ��"P��)��
�y��	�c�e�хI�J�Y��y���QĨ�J��43�e�ъ�=��O��~�ѩ0�IBա���@�@�P�<0�C!��8Ӵ!�0r��ЀRD�q��D{2&�r�P�;��O�_^�Qv�@��y Y,a�Lh�ؠden\����yB�U�2�C�iX`X������x�iNx�(Q�ԪP�1�C`@�p5��>y�'�R}��j�Kn�0@��G��%KÓ�ē5�����~YI��������d;6�}��!PdsI�b��E�3�\.I�����hO�>�1	 �p����ʚ��N�x�a2D�Z%mA<���Ec�u���c ���E{���\�d<:��$�%qp�y� ��!�\~�R'J��JT�cԦ<!��Rdbm��FC�^A(���B�!�D� &��59���XO"���A�)8!�� �Z�� �Q�8� �O)!�$��V���ʡG�=,��cOE�	!�$U�"�Z�!�A� y(B��m�+�'a|��V��mX��	� ��Qa�R4�0?�-O��ST�,��88�8H�
��"OZJ3su��sU�V�t�g��0$�,2ٴ�M�۴�Of�U2e�ԑ+!ƅQ�)B���'R��PK�0wxfK�"��m�H��1�4�MS�y��D�ȟVD��k�dU @�e�F���O��~·�8~X"8�aÆ.VJ�ڥH@y"�'���c&��*`�!��	x+̪>)L��(��Y��i�J&�9���~m
GN:D��C���"t���ԩ�'p����e2�I�~�O��˂?2p�`"�_T���' $��`�8x
,�S,��jl�<޴��'꠨�㉁��(	�N�(��l�eWSdC��#e٬][�N�h~�h��U�B䉷A�l��e�zVLaei�n��⟜�鉰n��A�x2THU&^�X�B�&7,`T�w�l�J�y��ij�'�M)tΉ5r�a�7�M61Dp�'�(�I�X�91�ɑ7��),H>�[�'%bаf�� �.��vK�:��p��OƢ=E��&�:Kw
ϝ]�
 �3*D��yr�ΆZ�>�wO�Y�9�ee���'m�zbiW�8\P��B�W@\L��/�y��R�*��
�2zB�t���7��*�S�Oav���?$8��B Ts�@�'&������:������/:����y��'��XB�EiRm��K��]o��
�'6��*�,X�� P`B��T���'Ax�oM�| �ɶ�A�TA4���d.�n�;p��$ܼ�;�KDu��Qi�"Ox���S��ϟ,.�~ez��b8��C ��-w���Gt�<Y��8D���Q�5$[�x��h��W�)D�(����V:��j����T�lK�):D��i���>������[bt@��B7D�� �t)�ȍ�F�!/S�D3���"O��mʀ*bfu����4j.��(%D� �pI78�ޅ1��t�cm&D�ȳ��O�>�z5ʀJŘXSF� �d%��ȟ����_�)7(E�KM�b�S!�x�'D��pN�:㞁��f�$%�j5�
���d�L����FL�D� x��T�!�$ƦC�&qb��@�(:�V�� �!�Dߋ{����6<��E<�!�ĉ�^�z���eN� N`��7�"f򜔆�@y@�� .�&u��|iv΂�.�,|��ȟ��OH���� beHT�dO��*t�ҝI��	��.�~�'���l��� �D�#s���'��l��] 5����╀e�Bh��4�~��'�����$ {�̍a�_��(�K���4&��?���MBx��˖� sbi�d++D�d����84�e[W�J6.���%j��O���ħ��/�v�Y圻��K�*��hƜB�	]袍cV��;����5�Z	dc��$�x#�'�ayb�����Fc��
V���w U���x2�ޟ.�H�3�E�Z���� �3x7(6mh�
���E�8��5��ǎ%nؾD2V,
�T��O*4���	A�uW�I2��:f��P k�j�!�ǕV�����F4$����I�!R��	�HOQ>��m���J�{lA�;���,5!� T���1��i�ܠ�M�*P4���>)'*B;F0ѡ�$�p�ڈ'�F�<�LU�Z_�H%	e��c���x�<��ϋ�I$t��cO�Kw|Yc�J�O�'1�O䠖O�h�O��j���X����h�)+	�'���A��"�b���*^�T�"Q0�Of����>�Ģ�f�!E4����֠i!�3C]pQX�N W>�i��a
�QP�_�l&��g�3�Ha�O���%:��тact�ȓ*$�(+t@2*K>�9�dܨa���ȓ5ю��@�4	�2�I��	�=�(i��c�����"���&���f�$�BI��%s����*Q�x�K���"5�^Q��:��Eɂ��0zGv�TK %�<��#f�i���
��TeM�kθ�ȓv� k�e�EB�䢔՘C�jy��)V����H�pE<-@�J�B�e��I�v� ƣ�
�=�b�8�Ʉȓ/�<ٙUn�
���u�K�XO�ȓd�S�+�{�	�c�%z��p�����e��Y��9&
�t]�I��P�� 1�(Y��Q���A?� �ȓ-��1Cdk��Z^�5�7�2u��Q�`=��NX$!#�$�&mC��Їȓ["4<����zO���&���M��V��U+S�0/bU@҃<7��p�ȓZG�ي&�^?�|��6>g���z<l	�V��$�Z �88Zh�ȓOS��r,ہf�ԣ1.�2fW�Ȇȓ.��-)��C�c�$8R�iäs"`}�ȓf�&<�b�
.^���c��%Jm���ȓ5�ڸ	g���K�����ʉ"6�P��ȓ5���GF�e��}����&Qv`L��:5�h+A��:��s���W{����qr0�Q@%yp-�P��o�&��ȓk�y#Re��.�ܬ`bG�5}�����}��)#ӡ� )E@�0��I�Go����\V�0Ň�e�Nܰ7dF�kԵ��%�܉����2�A䨂-&� ���S�? �Hg'��Jd ���3�=�G"O�a�#��//h��Rl�Y(܀�"ONbC�$�U�jN�J�kw"O����KP
M�`)$�Y;�"O�Qq�ʜ}P���g�T�ju�6�'�2�'Gr�'m"�'�r�'��'�048�̂#g�h�85
W�0>�d���'�"�'���'���'%��'��'r��g�<J���u��7�'>r�''��'���'���'�B�'�1eBϲ	;Z�jFk��(uڃ�'.R�'�R�'*��'��'�B�'a�a�T�I8*hⱺ&��4=�p�1�'�R�'$2�'�R�'}�'8r�'��Źw�P�mx"��Y�Lˢ�'��'w"�'/R�'ER�'�b�'���G�	S �]���+n�� #�'S��'>��'���'���'�R�'bP����F�n�fc7(�i���'l��'R��'���'2�'�"�'@���f��A�z��1� ���`�'_b�'�r�'�b�'���'���'"r�:�eć5����"xEC��'V�'R�'jB�'�R�'2�'���$e9
��	X���?.;r�Y&�'m��'���'���'���'1��'cB��.�t��1qs�ԧ%?����'�Z���':��'���'�R�'u��I�,t�+���b����ETjt�'s��'X2�'�'>�6��Oj�DX
)��X�B�?*"ts��
V��'��]�b>�b�Vk��=1�i�7�ڠ6 X�N��[�6p�Olmm�{��|Γ�?���Ϯ����@M�+v�̙�iĬ�?���<|�TX�4��Dc>=X�'���-[��`�F��%C�4PB�DL�N��b�T�	Xy��Sdp��� ��D��-�U��?o���4.��������y�O*
�"X�P��JǮcR杻t ��'��>�|䦅�Mc�'�La ˇ�&.$8ԧB6��	�'��d�ß`c�i>��	�٘$�1`�^m��s�»{#��	ByB�|�#a���{B�^Yj�{�J58R+��d����?y�Y�T����͓���7:}�����I>R�Җ�S0?���П��!��`�b>���'~����	�ƪزVJ�4�@���J�'��ޟ"~��L�:�Ć�%6�0I�hך�\�Γ+��ǆB�$P�Y�?�'*���p#n�� 7�Eɠ�m�.��?	��?Y1� ��M��O ��=��CC�G��0���!5x	)��H�6�Oz��|����?I���?q�u[�|�Tg@�?���B"�
xª �/O��lڶ!P�����h��]�s�@b�CÉK� ��?��rc�����֦��ٴYm�����O���� ��Ѐ��'P��@��]4?x��kV�ʅO�%���u���ڼf#��SV������X��a���<R�%`f)Ѷ,�a|r/g�rm���Ot0h��A�fJ0i��Ď�W��%�1i�OP%m�f������M[��i96M%bRX�0�ŽKbl��G��pИ��fpӌ��ß��g�K+�4a�Yy�OfW���Uh�"�#4�!3 ���y��'�Tᰶ�*J�J�sV��_��4��X���	$�M[te[G��!n�(�O6�Ȍ�zg�m:���^�z|*3&#���Oz�4�(\@�giӶ�p��$�
��C��}=H=ڳ�/���j�Ky��d�E�t4����z�p 'I?� �ٴĺ��)Ob���|r�$�
R�C�jZ�$>T5J�t~2*�>��?I>ͧ�?I��nd]Z���2;�� ��0P�L�@KZ;�Ms�S���S�Z���.�d��tʸ��D�p=6�Z�bn�C�'&�'��T*��Q��y�T�1ݴ}o
i	��T��L���]�IDQ�f�?��Z	���'��i>�	�O�ɷ(;=H"�_h�ٹ�o�"6l���O�%�""o���	��0z�@�:<:�i�<Au���"蠃���$�MSa���<�)O����O����O����O��'oz:��S�C;>�`��AL%d�@x��i��݂��ݣ3yB�'��dK[8	�b�'�6=�6����� D����0�L�S՘�;�`�O^��(�4�:���Oz�'�o��ɋb�x��"�3��0�T��9*�*扡_o�X1��O\�����<y�����d;�dh�*�> �� ��?���?Yu��d�¦���?�Iʟ���5$��ɳam�c"t��@Z�I�p��O,�D�O��OY�
G)6J�H�p�R��XD��<Y�>~����L��M��O����~��'���8��\ U5����W�8dne8�'��r�,_�SϮ1��m�C*Z�U�'��7�ߵU���d�O��n��Ӽ+�L��x����˕(a��
�C��<i��i��6��ئy�pI��A͓�?�2�J�_8��	L��0��ֳ7ԍ�6� "|e���J>�.O��D�Ol���OB��Or�8�˟bv�H�3H�)�����<�#�iL��0�Zk`R�'J���O'�'� �s�Q:eo��J�DL�}��1y�>y�������'��
M=��	�o��T�`��g�*��N"��	.<�ٺ��'D��'�Ȗ'�̈(�C�5��H2@O$`����
�J���.�b$�/aцPvkH�1�m�����yb�b�f�t�O����O��$N���@�g'0p��+��k:
y�Oy������4ruIG�>��i�<a��ο� ��`�M�|V e�1�H[���G5O���$��{�$��b��)���C)�U>Hʓ�?)�iI��ɟ�	nZx�I $<�x%��;�VQ#���2��$�P�IƟ��ɘSX0m��<Y� H���Wj�-�|IB<]�,�9c 'v�^�	@�Izy�Ă**y�e�^�p�j�
C/h5��h�4f�����?����ii��ȇ쓙�6=z��V��	���Y�m��4e.���4�O�R���獙b����A�
 Ln	(���ވ�塘\��	�?�bS�'op�'����eF�/Y�Lh������eE7�pP�4`�tA��Y4L�{�f��9a��� ŗ���Ϧ��?�V���	�e!Fx'F�q��#F �};X%�Iȟ�V��ئ��?)�F�@�2�Gy�C=��*�	։7��P��eF�y2]���	ߟT�I������ĕO�@��cș�l�&,+�'����4��	r�<۶��O����OZ�I��5~��wZ�����D	�e�1�Y�]H�j��'�O�)�O,��)��V�d͙64�X ��1��\" ��A�$���t(1��"�O|ʓ���W.,{,����O��Q�f!�Gaxr�p�ИK�h�<���$d�(�[<b�h�D����X��Ȼ>)��?�L>aFE~��3W���Bo�o.r�I��p�	Y��o��d��j�'��+M=C5r] C��"��6*�(0!��d] �GW��p��J+x�8��yL���%�r�'@7->�iލ� FA�r�-t�޼x��O�n��M���iJ(�R��iG���Od���&�*#T�\#��Y�KK�^���	�2v:-`v� M�j̀��[8�@ˣ&�lCV��E.�rU$�QD��&^J͠�F�Pj�!D��-Fl�E
�K=���'x�☱��ƳQ�h0XB�
do���Ʈ�O��� �_� 7�ɗt�T��wd�.1���2��6D��T��/{W4���b��#�$�4NK{�@�6���س��<P���m��氁�`��<t�0{���I�|��� rc.�� &	�] ��:�e�2�V�@ve��\�;D��	q��A��-'�l��/�R0H��Ƹ	�� /)�2DM�;G��5Cܴ�?i���?�����	�@��EQA*H��4�7��_	7Ϳ<Yf�^}���O�m��K�����"�8p��شT�h�V�i���'���O,O�����K�8���$8���{6�D&޶l�yU"<E���'/ڈpk
	O�����*f$%�s�|�Z�d�O���h>�'�8�	����1��]�$]�k]�a�c��8����>ѐ� `��?i��?�w�%�4�p��$� X�$�҅>%���'E6d�H2�d�O��$4���zD�0N�ry\(��ր|[L�(�P���g+�I͟d�I����'�~��/Y�@�-�4��#?�Y�E@�T2�Ov���O$�Otʓ�敻�nQǚ�pEZ's��̂*��I�1O����OZ�$�<� ͪT��IƜ� ��[Ĉ�J#(��O���QN<����䓸�>Wl�	�T�N�b���X��X��� ���?Y���?!-O� Ȳ��{⓸O���AH�\Qh��&�Ҥzg^�ܴ�?!���$�<!��N��OJ)j��֬)���3�@8`�HĈ��i���'~剔< �QI|��j�b��B��� E�L��& �@��'��	�,�^"<�O�r��7@�<GN�pY�M�%#��kش��\�!�=��'�?���"J�	 �x�q� �A
Qg�G,g��7m�<��|���OJm�%�+y���ɰ��� �6E0�4����io2�'��O��c���GC�z�8�W�ۙ5מ����M����W����K�Y>^m���u`�H��(�=~f$m�����П�)���>���?)���~b���$�h�A4���"��_���'�d�S�y"�'���'���P�ōI �,�&톖T�Fhpac�L��L�4�$���	۟�$��X�J����Į�Q�,P�SJ�2J�%P�<���?���?��O� xi�k� "����%.��I����O��d�O^�O��D�O�pHFE�1K$�Qt�ш��#��Q�a<:�G����I�����ğ<�ɱXl5�',4�!@�9u���s��R̤l�gyr�'��'�b�'��y ��ڴ�MK�F�&��y��!�.���L|}��'�'g��'��-�0�'"�'	6#��1m|�{���&7R�9��O{�@��-��OB��D&�T:tl�+��!Z0ɛ�l��y�fm�,���O$���O�xШ�O����O���럮��*�c�����9rl~��f �{�۟��'^j�������F�:j�Ad�`�r�෿i��	�SY�<�	��	ܟ��kyZc2B�
⬖���9���2xDL��4�?9�(<K���IH,oZ��37�ً|�^�`�n@�M����?���?����J/Ob��O y���<0Lu&�N�]j�h#7�����0���h�S�O�r�]#o��͒eL�9%�����X��7��O����O>����<9���?����~b$@�J,�I�W*�a�E�H��M�N>SbR�X�OLR�'�¥ңh����b$�1�R�����}/�7M�Od�:�F�<Q��?�����Ӷ��3%|f�)��U�Sp���o}2�!E��'���'�r_�@{T�r�vi���*~�h�3�ğ?�D�'��'��|�'�R��3V���X-����&�;��X��'����,�Iğ�'F.���П� b�PHҳV�Fm� �����SC�i��'��|��'��)@lm�d8KJx��J�� �XA�A�=h��I����ןD�'��U##P>U�Ƀ%���ʙ�{QA����pH��Z۴�?qI>���?�挀1�'�6��Sc�	\���2DH
.nc$Q�۴�?����ҍ6^�'�?���b��E��"��c��08��U��FsW�'q��'�����T?I2*��`'
�&6���ak�D�s�(����?1��?��'���P�#��E���P�wB���`� �ib�'��$É��)���<���S�/�E�W/�0���W�"���'���'���Y���Iϟ$�����\\�c_�|��ea���Ms��A��������U����,Y6_2�Qx�I��O��Ul�ǟ �����C� S ���|:���?� �)D����O��*�IJK����'"�Y���������ɍ
�Tl��d߻H̾��ҮI=P����4�?Y��K5&_�����'OɧuGjE� �6�����[�L�����?9/O����O��ļ<	�#Zl&�0�1�,pzT����u!���Q�x2�'�"�'0�̟����Hg&$`�&�]��p;��[�iZR�
�ɟT�'���'	�I���yT�a�s��[	H���
.�m����ʦ���˟��?y���?��U�Y��oڕ�ҝ��,��
q�J�*9�5�x��'��	����O^P��'�ұ��KE�?�,�S�ă�M�׎}��㟰�	���@��p��O�h�C&��\`�a�a��=y�iA�R��Ɉ6� ��Ob�'��\c��p�] x��i *�Y��ZI<����?q� �PD�<�O�0�p���0N�$��Ӂi ���ش��d�9�dAo������O��I�t~ҏм
�\�pM^i��}Â�ۓ�M����?!B+�?����O��s��}��R�:R�B���{N���`�i��%8�'���'B�O�)����A_��2'� 8���c!X<F�v*J�R�9�y���O�}ჃH+�L1�t���4�qa�����韰�I�y�:��M<�'�?	�?���@w�8r��=�ʞ%�p͑��i�R�'�R�P0'�T�g~b�'��j���P��l$<��bꁩC��6M�O�E�2�Yg�i>��󟜖'��gD7 ���#C߾(�RE��fӎ�D�#2b8��<�'�?�*O �D�-2�����'���c2@^! �`(��n�<����?��B�'p'�+q�X��CdP2U���!&�O��5f�Ø'�rR����'�(����P�ђ$C_&�AP�����9m�̟���T���?��,��-R�YƦ�A�.PvI��Cϑ5e�����(�D�OBʓ�?�vnI���	�OZ�I� p!B0+�?�"�Xs"Φ��?A��?����g�i%�`�1f?l��dj��'�EI&�p�j�$�ON˓���X��t�'��\c�Z�c�Ŕ4�.!hg� �^Z��۴��$�Oz�DH�J��/���kL��TL����G�v������̟9$�\��P�	˟����?���u׮.7�E��>d�\లA���M���?YdHՇc����<�~0!B#v���K�G�D!�����u�V�]�L�	���I�?і��	B�<�rM��C�6�d|�$�V�\�@�nZ�x|N��'�)�)�'�?�4��8?H�C��=n��P4���5D"�O����O\4pD��_�i>��������)�'M�u�����0�Z#��M���?Y�d��Q� X?�	�<�	ҟxҴ�ç K�Xӵ!Z�)��%Є��M��9�m��x�O3��'剧 �5���/S�9��ZN8a�4�?����$�?y+O����O��ĭ<�S�	�gt&(( NX99n 
ЊYM[`�qW���'�BR���	�����?F�
q��L&5	PmH4�IP)P����{�D��Ɵ<�I���	dy"�U����9�K�y��)�!�=(`�6M�<�����d�Op�d�OX��gU?��� 9~��58#�Q�X��+f�f���O���O`�7�Q�X?�����<i�.U�G-F���6u�ԕ�ش�?,O����Ot��ߖJZ�d�<�!�5^����N�{�c��ԗ#���'{�S���������O����X���kSh�����jx�CfOJ}�'�B�'i�@Ο�ItJ��_�3�F98p�<m~t䲐O�Ʀ��'�X��3IwӤ���OD�$���֧u�+I7&h4I�#�q��A��β�M���?aoJ�<I�Q?��_ܧ<�> �@��{B��@�.���l�$O`��ٴ�?9��?1��*7��kyr�t��TC>�>41Do���6M�.��0��.�����cf�v.|$0���,

b��P��M+���?��*��5J��iDr�'�R�'�Zw�8�p��q���WAӖ+����4�?�/O�T!�2O�ӟ@�	����N�>eW
ll�A'M�
�M��V�jvQ���'w�]���i��a�+D�%+�Kc��&|Ѽi`��>�Q�G�<����?9��?����D�?l����4�F���1�(`�L�*U+Ez}b_���Nyr�'pb�'�T�����E�LI��@��BH�A��3�y�\���	П4��sy"�߻�8��h�D�[=�@��m�j�Չ���'�bZ���IΟ��I�h�i����� Ҙ:��.XL���GpӤ��OX���O��d�Oz���(���5�I۟l��!��]����V�Q�B�8�f@��M����?�����D�O�� B�7�ɞ9�@`CA7�Z(JJZ�)��g����O
�d�Oh�!p#�צU��ß �	�?��
� �\)��ݲlD��*��A�?u ��E�ibR���	�DT��SH�i>7�T�k|n$���ߴ��X{�d�w��f�'r���n�6��O��D�O���������~\�#�7��<��@A��' b)�#3�'=�X>M��x�"�ì]����W�~�P��i�$��%������OB���4��'��	&,�ypH��JF���5����Ubش}�y̓�?!*O��?��	���q����i����+����4�?a���?��Ί�@��6�'�B�'?��uw��A�,��#���[׮�!�MK��?��P���S���'�r�'q��!	 <�!��f��r An�6�S�Ά��'�I��@�'Zc;ֈ��:v�⅏��T�P�OV��':OB˓�?����?-O,,Ȓ�D� 		E��T9�X8�c�7����'B�؟4�'C��'c¨ƶQ�U����|�p0�Ü96F�қ'��֟���ؖ'׆9��t>���T�.�<<�FI�i� ���lf� ʓ�?!/O"���O���̖U���)7���A�M[�6L	d
ּ2��lݟ��	ğ���Uy��΄ꧯ?�c�G�(P����.�����X��f�'��Iϟ���џp�iw���	K?�E/ύ�H@� ���d�8�f�A��1��ٟ��'�n0���~j���?���47��#���8YX@� ��o�0��R���I�x�	Z����]�W�e��&e����G�xG�}ʁ����ٗ'�v9j��s����O����&}֧u�g�:Y,���k�~�h4�MK���?! o��<��]?���Y�'x醥��m��Ks'V�b�P�n��;E�aAڴ�?����?��'PK�Ily�/U�-=^e�g�ڜ��$���x=|7�S)#���<����O2�8G)�ة�B+
��C".��DB~7�O�D�Ol<�1Ho}X�\�Ij?Q�AM�+2�t!�"I �[c�r}�Q���.?�'�?Q���?Y���u`�J��	�bq6�r�	�����'��Ȱ�C�>�(O8�ĥ<���릇��U�<�@�,z.T�`��L}����y2�'���'�R>�	4&��@�曆X*,���a�2Ƕ��`�:���<�������O����O �Z�H���xҡ�NR�r���
b��d�<���?����07#���'D<H���ҿ6�XH��I1V
�'�"�']�'�2�'���B�'
�y��.���Q�F�
&���p��>����?�����Lژm&>��D�ܺ8׾�٥,X3���0M��MS����?Y�h��IΓ��kD]B���b�c�D"u�նiw�'�I�Af��rL|������(Ȧ/6��*r��g,��2SηQ�'�r�'�b��'Cɧ���v~R�x7��=1����C9(A��^����E]��M�T?����?u�O����8Wݪ}Q�ϟ�~>P���iC��'������'pɧ�O�����ǂW:��f��}��ش71�q0պi�2�'2�O^\O��Dܷ^���[u��Wp�z�Q�m�D�o�� r�?���t�'���'W�+�(EB��ΰ_5<p!��'yr�'L�4W��O���O��I@I
�3�#��8����X�7�)����.��?�������	�B�&t@G
=$׸�ϑ%i��4�?�`j�V�O��d"���x9���F)�"�13$��Wɜ�pQ��Ӕ�j���'�b�'?�Z�P��1��@�ポ�{.��
��`K<Y���?AN>Q��?��o	;���E�@.�l����(�y����O$��Oz˓V��˵0��D1�OW���u�D�]����_�p�����&�t�����ڥ�}���͆o]|��B�ʹM�4(�-���d�O����O�ʓ0��}y���Ǜ�;�.�����F&j)�׌$L�X7��O�O����OZ�����O��'��+�!��~J�%��a�4d/�q��4�?������F�6$>E���?�+���v( x��ͽ�^e1V����?����l����S��c��n�[S�^�cp�q�
�M�(O��Ig�^Ӧ0�������8�'$X+"��\^R,��I��+|(�ڴ�?q�]��D���S�Qy���.�"�(ђQH�;xBf�n�
q���������	�?�aM<���$�,�(��$"H�;DE�=�\���ib.�*T�'�ɧ�,�d�27�d��eI֦3�0�/�|�^@n���IӟX�ݵ�ē�?!���~�ȪE���E�ݣ��*#�2�McM>A�O�"e�O�"�'��jQ�2�����_�X\iz
H�N�$6�O򀳱�_k��?aO>�1>�f鈄��A��XG�VQ8	�'ɦW
]�	����֟Ж'�J�J��2	.\�:Bѩ=z8؂E C��b���I~��ޟ����j�R�r�jEU���/�p�,d7�w�x�' ��'��Q���7�C���Th^�*<�.��I�| �ɞ8���\6m�O0�O��D�O�)�(�OdT���I!�XH3���b��
�O�j}b�'�'���'� ��q����O�ԱG!��l�y��gp��Y�a�����qy��'��b�O���O\�jtⅼ.�@:#�O�PyxE�e�i�B�'f�'<PM�U�dӸ���OP�����	N�I8# �zd��+d���`�m����'m�Ȅ����'��i>7T?B��۲dG0 h��[iC�v�'?r��ܘ6M�O���O&��䟖�$�t�(q$���F� ]2f�"|2�'M�*�*��'S2\>���ThiFědOpA�@.�>/�tHr�i�ft)C�i����O����	�O@��O,�� T��ƕ� cx\"�n�A#�x��i;Ty��'bɧ���d�'��8��C�D팑�D� :P�T�`�lӂ���O~��^
u��m�L�I�T�����]����s4E�z%ȉ@PCF�ZL7��O���)����?��|�)[��:G������Qy�E�i���W ��7m�O�D�O����D�O��(f��:qFDP��;n�Hc�U�`h��g�������Ißd�I\y�)�� H�c�y�3�K�[��T��î>�+O����<����?a��\(�#b���3h�!�u�؇;i8t����<q��?���?�����ǎ1W��lZkp~ 9T��V#��[R��!�М;ܴ�?����?���?*O�dL`C��ȡtU�4�0l�K}V̐##F�K�ޔmҟ��	ߟ0��[y�Ѻ;�`�'�?I��Ձk�<�1W��'�=�sEIV�f�'���ݟ����`
u�#?�禱�X�q3��*�ɛ#J�x���kc�����O:�#I�Pv\?Y�������bx��be���T/��8&U�	m�T�O����O���X�*��$�O\����B\D��hE��7pֺl��͏��M�)O��Xu�֦��	̟����?qڪO�.�P�L�����/m $�>W���'����y��|��I�
i*St�-=fƬ�pm�3*�����e:h7��O2���O��I�m}Q��HcM�`$�s���SB�q;�(E��MK��<���d-����0�(١�A5P�W]ą�1�D�M���?����|��7S�@�'T"�O&��t"U�+�6���Ϙ�
�:��@�i��'���X�����O����O<��q���<���H
�#:��jR��Ħ��ɟ{���O,��?�-O.�����K�c�<�p+̚l�l�ix"���y�'a2�'���'��I^6<AJ
Bi zI�/�
Sհ�ѐ���$�<������OV�d�OjeRc�*_#���@��]�
`��G[�9*�$�O���O���O�˓`�JБ�0���85�6X���*c/�a�2U�i��	����'��''�����`��ҁ����������4��6�' ��'4�V���5�̶��i�O�ze�'_("�a"Y�Rh��'�F�E��@yR�'4�'(�X��Ol�ia5O�F�zT{WGۆO ��f�|�H�d�O��<�z-ېU?���ӟp��8-�}��-Υrή�*1M%~��%ѮO,�D�O*�DI.|��D2�?)��ɒ��Љ��)ǄL�x2�jx�<�2k�L�i�R�'��O��Ӻ��Ϟ�)N�q�gAC-�Zt��aX�������Q�|�'�d�}�gk���HM`w�Y�&��@�W�覕B@%��Mc��?I���7Q���'`�$j�t����玉v/~ap�gf�H8��9O����O��d4��П�d@��2�Տλ5|Py(o��M���?q�]��c�Q��'���O��G,D_y��)1�ٙve�� "�i��[���dem��?�����LK"��&ᖆ`�D�s%��M�+���'\���'7_���i�u���ͳl�H`���6)�X�cd�>���]��?y��?A)O4𰴮�.v&�$��ό@�|�8C��t�Z��'m�	՟��'l��'Ur���e�@�P�վ@2c��,��|��O���O��D�OʓDl�YS7���:���>=�����+x3��s�i��I埌�'���'��O͛�y�Nɜ"i`@`U��b?.$���]����?9���?�,O�@+��E��'h`H�v ��}��0��� �;��y�үu�����<���?9�*$�̓�?��z���oK4}z�@8q���Ӱi���'&�	�i�dԙ��\���OH��<
<�)�M1`>�;6�	 J:���'��'O�C�.�ybQ>��p��c��YO �c�[/2�ʁ�P#�˦	�'P�d�Ue|��D�O"���Z�קu���;-��H�g�Y(+D�@7�*�Ms���?�'Ou~�^�h�}��f�-�N�����tL)+e �ŦY��������蟨���?E�'���[��@Q�[�,��MR��C�n�~i�Ot�r#�)�ޟ�Q�&Ƿ!� r�E &f[�e3Q �5�M3���?���n�8�rq�x�O���'��l�@V�&����i;E�� ��"��'[5"b�d�����I Y7��ᮚ�@��ʵ+�&'�Aٴ�?q��� ��DJ���'��'�ld�T��EbvE������$���g�������I۟��'��A��GM�8�aEŅ�(��`����+X�vb���Iퟤ�'��3O��8QcƠ>lܳ��^�GH�hH ƚ3��'5��ِ�/E���E�x��ȳ��ϙ��	I�4�v��E�ۧ�Z��3DE �!�d�N2:��DY|�Ĵ@��*#�qO(0V�Րgl@P�aA= �b�k'Oiaf}�� Gp��B�[�Oo̬[�m�4;u`�Y����&���4GοɎ�Ґ�Ȁo�y���V�{<L�Sj�*�|6����|��!Ί�w�*u�cAI��Y�"MU������S<n����	��!��M�A�ȡ1 ��3v�-!�'$j��o*�I@��,�6�s@�'���QN��ps��O�!U���B��USf�����3/v��:��l����K/j�R0d��ǌm�� �Îb��vcj�I�;��ӎ7t�Z��3
�	�"I��t��'�+��?I����OНy7e�w�F��A͐�a�4l�@"OZ�˅dځ $=!fF�n>&��',�#=qւ��: TY`�AA��@��e,�f�'5��'p�б���'��'���y�o��b�\�S򥈃'�h��sƗ=��)A
Xa}"���>=���L>��B��Щ�� QR�(�����<+��c*�>�UO��0l��>�O� �p U/�
W��1C��<��y�7�O�D�Oh$��/�Oq��	П�rb	T��T�����:��oh<�e�VHx��v�A�����
\~=ғ��<QGJI �Q3��w��H��,џB���A���?��?�����n�O^��e>ei�芃�<=�ԁ���6��_�jB�I�'�zx����
VR��-��0L~���+�|��f��&�z��V�"?��p����<ɂ�$�Ox���O������P�I�	�a�=l��	q-�"�!�DC,bPĠx$c�+2�<��iڢx�1O��'�削U�$��O �䕗__LqA0aϷ��Gh�(,� ���O	�� �O��|>18s�\�+l}��LQ���l�nIq����Iy��+��77ѐ����s�]`'h� ���MsH2L�ɢ%]	$�|-#�l8��)1��O��$�<Ѧ-ݣ%@�Y�O��)8�) ��Gj̓��=�1,ϲ	�6]I��о:���K�
<Ƴi�H�b�Ö�4�v��c%w�8�' �I�e�N��O8���|��G;�?����f�dT��WEh"��4�?a��IU49��̈Ċlj�G�a�*���'f�jњ��{��X�5� �ͦO�E���d.�ۗ�W�n�"}�� ��	�2�S ��|�> C.�B��8���'a�>A���x�r$CchP R�T�eg6�C�	E�h+t��L���
w�3U?���^�'b�db�jW:5>x �0t���2Fl�P���O��Ĉ�5B��g�O@��O��4��͸%g�+����΍� ���%>�	)c����'�b���$�xFd��CC�
��I3�{�K�k�nх�	�k�^���U �G�\�>�����\~φ9�?�}�����I�d���kjX�;�*�`�w~�U�ƓLW��kۙv�~e���D�?o���'�"=�O8��,�J왖! !�C$fX=NL!RH�)e"����0��ԟ�^w:b�'���B��ݲƀ�>"�F���+��	c\�!��%Jc6���ܿ}�$T��/B�m����)�1cB���L?�̤����[�@��?f\���-�X����]�!h�b�'R�'��V����v��P��퐍y^�ٱGI���x�V"OЁq0�U�GSF-{�KǝSľ��b}"V���$��M���?��,� :�aqIS�6/��zA�ƴ�?!�B�
��?)�O���@�'ԤIظ3H�)&��J��5_����o�(v����"��t8����@֦m�3w�Ƒ�@m2g�ӌB����č'�&��B�5B��x�g[��?���?���R�Ȝi!M�9�e�K�c���j-O���%�)§�r���Z�^3�][-��r�Ն�dK�&k-��=��̏^��@F�Ͻ�yr[��������O�ʧ0a6��!�̉���YB�a�`�,�������?%�قr`����	�>Of̑��"bg�}q曟��i4U-V0�����anJ'O�('�~*xiwHZbn�H�R�ؤ�Q'H�v��'X'���eʥZ��pתC�L
ŧO>䃑�'�"�ퟠ�i�n�,P�g��\�Έ1� 1D�|HQ�E8��}�����L�E�$O<Gz"ˎ�FEĤq��58���^�	����?a�"�40�/ӡ�?���?��Ӽ�b	5M ʖHJc�~�(6"ϡZG�p�7�L�[��˛�[F�Ҏ�L>1eާ'Ą�Y'AZI+��P2�d�]SQ�U�Bu�G�FP1�}&�����L����L��[o�;bC
՟��	˟|��L��>˓�?)�G�,g� �E�G�>�G��9��x���ls�1��,?�ղ"M�����M�'I�UyB�Ěmt�@�OݩH1��!ч�:e����g�Q��'R�'iv�'�?A�O���%.�NxT�Y3"��_֢-�U�\	d��B�,��M�Pǐ�ul$��M�oߠ`�Ο,<LiĤ8f2����?Y��!r�F�]�.�зND e,}#g�'�2�'��V����W��\�R��)� �1�KQ�}
*��ȓ8�8�T��,*�ĉ!���l���<QZ��'�@��/tӰ�$�O���lJ8t@B ��ٱ|�^��j�O����[��D�O�S�D'��˲�U�l�����'�6T��%�]���I"H�0Mw�l�	Ǔj&��� I;F�Y���O����N��B����^�P���p<�D���$�I���I���R�_��@h��]�N��9
V��<9�����*x��K��8�btrt/�/�>Xp2OԅnZ%^�!�dܑ-z�M9�i�$1>�Fy�G�6�O��ī|uEK%�?2��"�qa���c�5��,�#�?)�~��pb�'՟��[!n]�%t*�jʧ*�� ���@8�{����1����O��D�\(8c�y;C̄6v.#}b���~�4]�%[8/Hd��d�Y�ʶpQ2�'R�O �π  1�A�&9\Erqlڤ\�����$�O���dF;\/l�	dOM2�4b$�ъ4Hax�l2�RS*p4FV >��K���6��%�i���'�" ��!x��r0�'p��'�w���q���CCT����2/y� (�9.��ɯ^0Ƙc%c>�3�$�:�(�3���7��Rx��@�@����3�,� �C%�3��\�om��4��"��}���m�p�mڷ�Mk��g�6A��S�gy��'�jlX6�ڇt�j-�d�>k&�[dO��<1a`��`��w�^�xw��<ۈ���~BR�00'�\�n��	ӳK�:|�t!k@������+�������	��	�O��Su���2�W�$���ោ-�.}{g�h��̋��=��m��B�{�(p�&u�y��ɇ=��I0�T�j���S�5J��\�^���'EB�'L�ǟ��?a��ߛe��i��OYˆ@ �`�k�<��*���A~iJE�c`�`�	���hy򊂟.7��O���M+1���dUR*Z��∘��D�ON�x"�O���d>��CH�P ���ŀ%g�(oZ$���+&ʉ�Q�b)ۥ,,$m ����0F�T����R��om��mb��1��Daf�� ""�3B�'�¼K��?�(O
�a�X�8�� `����>O|���O��"|�+ʼ=�hB0,R*8�8H;J|<�i�����E�J9hdH1����'�ў"~Җ猀w� �#ÞT��ݡ�� x�<1�ԋDx��*�
�%i2lI��p�<iፒ�p!��"'˕ukdm3D�i�<��k�7 �SUƘ�<1�B�Jg�<����+Ȏ<�Щ��t������^�<a�M�[?JH��X<��7m�T�<��䏋sW��!Ꚃ#ʨ�q!�P�<�p�C�|�\q3�Ԁ@�R͈G$Ht�<3��0eAs�%�9R+N�Y�u�<	��~J�pK��J�xk�Iy� t�<y���2i��l�B������^q�<���(e����4��P8U�E�<���9��`��F�8��,�B�<y'E6�@�Y�hJ�+&��3#�}�<9�(Cc�L$C�ʅ��HhUd�z�<Y��ؖ8k���͓/����u�<��ھp�X7��h;�)�'
U|�<Y��	��m���G	2�k��^P�<�V�  �JL�I	Yht�e�M�<ٰ�XU�0�2N�9F��ŢQ�M�<�q
D)z��HP��^�[iRH��a�<���ߗ;f��yAdW�R��`_\�<)�%��PvB���.��Wp�i��*\�<���to&HY�P��P!���\B�<��'��88<�a���*	Ʈ]3�Q}�<��	^�Ur��V�/;��}��+�A�<A@h��U��]yr���Z��u�<�H�d|
)����jw���D�Tm�<�W)ۡU*j]AE��n��)yp��;�X���5�� �I��Gǈ@�}�H<Eg��	�m-@��t��_< U9%������it�H���� @:�9QVi\�0�ع�BϞ9k(	 �k)O�}1��;x"�qX��F�Z[(<q�l�7#H`��#*�U�nu����3�p<��8KN�tb�j�X�r��˝�Y����,[V*�i��ɫ<Tr����d�ڬ����(�~����<�r�*��6ل�0��$q�� �&lO&�� &�;D���JQ�N��Ȱ!�Ҙ"���bҨO�;����/�::��'FuI�O�*�+���f�u�7�[�x��r�I�D�u����0$lb�`�B�X�����TZ��-�"/B��'��*�c��:��%H��p8l��剎�F7����Y� � ��F���hpk��~H��?Y�#��gOV�'�(O\$1 Hߤ�R�y�l��=2|����U2C�'st�B�阩`��ۜ'��V�C3?lq �̄��%�V�\0-�<3���6G����ėbU2e��K(!n�ԈȺ6T|�'�Bҩ �1��rì+ڧjsru��B�M{xS���O�$�!��^}� B�:r�rt0�#���rjȃ��y`�4+�!sV`ڲ����#��ӷ�:� �#o�a�1r��Გ� �mbp0�5��5�65Ey�fB16d���q��D�ʺ2��a�'� ����NԌeMXe��GZZ�¹�!�>O`T�R�D�o�Ԣ�&�;^2��� NՎaEHE��{@ΒB�ҌFmY-u:y��d��k #��y���~���BH޲8ҍ�eHq2Y�3�*�yBd�u���J0E�:.^v�J��TO�F�S���D����mK�����	�7�^EJD�X�X�*�y�"�	{z�:��T�@��ʑ�S��r��#8?i#FE��$
�e�1mR /����z5�|�O�3���̓�|�	���d����]Wr]H�I݅*�\�'����,��iZQ,S,Ԟ���C�H�>p�5�ce�bp �J��e�+�HOL٢`k��<9�^G��A�6ƅN>&}jv�1!�e�w
A<3��#�b���R��O$?/ �1�Ѐ���*�
5)�E��
0�I�~)� ��'�;E?t��c��&i\c���k��f�\T�J�~���pK�+e��X(�d��Y��9��=��B����P�CԹuʜe��
��j��'������Z�y&~�S��]��hB �?)���c��q}���q��$P	����O�@1�S>Iki ���Um�"�֘����Q�<q��ӆ^X��҃�D&#���d�.�p<�GC�S��!�G��p؄��3yj\Lc$J�!p]d��a	���=1 ��,[�,�D'r�$�&B�<���f
�3���R��>9u��4����H�<�4�|2-,pR�hC���(�L�y�.��O>n� *O��0��m�T}�uC1iδ �c����O<ɗ�CҘ�sp%ŗaޤ���-س<��ї'߆�OHa��ѵԸ'|"�b!o�1/0.� �Β�.�8�	�/�Vr���<���w�2�s@D�#O�����/�85RP�On��O���O)��i�#*:�5(g쓔��w���R/����'��r0o �s�ʓF� y%�ǥi��а'��5-vz ����a�.L�A����h���� ���.!N�V	�!/�\�2���5c� �@,O�!p�Ü�OW��' ��O�	�N��� ?h5l`-X�U�2��N�P�R��6@V�TZQ�������'��Y�獄 ':t
��Œ�B�k4�nӼ���'A4�ZN�擮@qO���5��?|����
�[ܪ,�Gj)�����	M,�8�ǩ�r�����sf��|��dF	�❢ �>M&rA��B�DF<L倌�¸�MB6���a%6Yb��_�{|�yK�J-Ld:�Tf;?��'XHu�/�*��G�O�����'�E��*�v0�B���}y���G�	bL"�q�W.{b��W�ڞ|����On�� ���{�.ʂ4$8�1�.�h2�����gi�-�7�`D�I42Z�ҧ�t�Ә��x%'�c�45�Ǥ���MwꅞQ/�e�f���Fq�U����ǟ�I^�Ozhi�QU?9A�l�Ls�ɪ����W��y����?����O�4�4[�{�b��j>"�v'�!�����?�y��+�O�ULX�Y���n�����Z̕O��0˃��t�,9�q�՟N�b�`���XpT�Ћ��A�M�vL��_!Ʃ�B! �D#���T�����D��OH!�C#�øO�٣������if�ֲ3&�������ArIVu�'K͚ �J�+�HM��U���@4c},p��H��Q��a����@0��
7�T(�O@H�d��O��R4�C3Ҁ��۟����k�Lě�႒+t2�CsX�\yb*ΤL��\��	��섁�
څ�rl�vM�%Z�@�:�'IN�)gJ�+�¡�S�J�k{<�B��"�ź�|e�U����d�N��'aP�tR���)rɓvG�7;�v�UF�a%hy
�*�	7T\��l� ;%�tT�~�ȑrG�{v����-��̎��xs@�&o)��)ˢ^O�y�T�G��i�
��ywl_)p�qY�n଺��ǽQvD� #��~c݇`�~�9�':�i������'ҺX�eΆ.`��t떉�9(-�[#O:Y���C���c�\�rW��zË�	~z"�ٍ�L�(q��M?�� �3�?�b�O���g
�?��F	� '��A���!7�IV�9�;AȊ%��U
x�9��I89掸��P�*�d"�
h@2ɋ�5��<i�BόmO�'��ɖg�8{SH�	�̬�=�%�$��jp�ԁ}fd��̏>��CV�P�f���aJ�P�|��)u��ht�ġ=�d���3֫I0O�	���<r�7o
*�MK�Y{����O_��p=i5mS)���H�.�2p5�a;v�߄v���3"�s�Z�Z��%L���J?�����Rjۤ��)��mHvb�s�I�
.S1�G1��� K�iK	`�C�'a����G��,:�16���0���TP�}0�)Ƞ�>�%��2�p��I�sFf�R��[� h'E��]QR����I�M��՘'�K�E��Ҥ��'��%E�x��7EH�DT�D�]�(�ɑ��T��xS�ӧ[Ҩx:��\�(�
E��0|�!���SI(�o')�����Q��ͺ0 ��k ✸K�z !�ʌK#@����f�N���[��Aئb~��O��u� H��vk�ѵ%��4�&䩰�I'I �y�	YS��� �:�oƙ#< Q�@�;�b���HyyB�
!8dn������'�n���Ϗ@%P��2��25��C�Jȫy���)$�'���c!�Ŝ,�����J,T["��6@iHmh��2$(0��J����pRd��"϶ HGbSe�� �D���p� �u�L���K����"�2�	/���&��+��AYc�\1|��c�� ���<}�~�����Ƭ�R4��O��ѓ���N��e�J#�"��I![Ԅ
B��$Ka8��]M���qH]�`�I����^{���҄`-�5�uO>�@�^(e[ L
�*O#�0=�B'���ywc�X�
�OG�<�ϊ��?��H1V�{��U;dl��#b�|�N�:u�ɉ+�<K�vd���O$'V�qx\y���=9Ǯ�Aѹ( ��υ.@��%��[Ǵ��;r�@�H
�DEߟ� T������%i�J��U3��i�� kS�y<$�U�F�*�ة����ot�hp�V�jir� 8�BI֩BO�G��тw����3�2*�j�A�L�Q��Ոc
�gUN(�V��8�p<�R+�	\�T;�'�ǪS?y0�l�N�� o�YD��1,:�у�ڄ��O�z'��¼CP�ʻ�aC�=1d�8Qu��{�g*�<1"�O�3�*Y{#nA�7Լ���^�8���i�M]+�HOZ�ڢh�:�{E�ŝJ�<���*�Z}���
B2d��ؓ�DY��H!�(���J'a�����Y����xt�v�Q�VI ��h�FA!�Q���)���"M_(��%�ѣy
4p�(� ��OP� 6``�J��B�B5ā4�i$������i�Q*P��0��]w�� a���8c����ϓ$]A^R��"�.�1�C�ɟH����G��B���eD�h��ܲa���6��LA�$��F���b�o�'���alz�$���AK�Io,��NO�\��O,�IS�굑W,և(�R-R�[�T�0�i��6��8�2����HO���%#/*j�ʰFT;��@���3עW�b��D� �ޏ+Ϡ��}���h��Æ�L�͊$ Œ����0Sv�
��$�83Rj|�` ���s�
��8��+1�l�S�'���0mG� �>����KKz��%J��F�$x���C���,��
"yj D�7���l�E�'7Е��GH0%����D�(�<e���d�-4%t��O�	�������GAȠ��/�.* 3�����^$Yaz��W;��hA��9�0U.!��3�h���"v��**2��q&`�O�J�7͘�X.����'6�rf��*��A�C�Cax�)�;p[��OZ9Jt�Š9�8�h�#�B�rLSN $,H-�s��f�b�#� �$qU�@ƂՀy/8�=	�c��\��y(S� �G��L?)`�S�,8��z7f��ݴ�(O�Ҭ�"U�~�9!���A@��B��mM�(1��W�(y��.d��C$�R�^u*���tb��pE�[R�X̓J͢�8�����D4�ԙ�H��J�#�c�O����5� ���8�
O�5�r� ��� ؐ1�$c� ��<Yg�A W�2�Z�M9�:�ߑp��e0�n��#�BG �[T8">9�C�L&��vh�h��r������̹<�@18��
9O#�<�q$}r��52F�{���b�>�;����'?L��*�84s���"煄h���'*B�A7��o�^I���A�?�L���D�jT������v��,����7Ĵx�B�8� �h#��b؞`R�c?N���d�0p2�ED5����d/�OY{D�H#g�&��KV�q#ֹ8"�8�O�� b��c���K��-���@�&72b�
ϓm��B�.r��
�&�1/2E�c,�(4VI{tJ��cfR�s�G+�<8���s��8`�!�<2�B���'��\���L�t��($����D�04+�)"%�
�"!J�5��!�bY8B�_:�6�q��[�8��b��s��K�x ��U"��c$�T��c#� f�r}�T*�U����\�C+�b� �%��Za���Q)�z��&�2�*�b[�L�&e�.7}\�b#����J���
��<a���
04i�3M�0?�lB$$�yҎҟb���J��ϲ~l������<I��ߒ>�����=Fm(�+��ׯMҐ�r��6V�p���0=�E�_;k�@9��b&]?~l �@�,|kT��..t2�0��^�	P�2�2��>�d���N�?l�p�у�yN�)ԁ��Pd�8��)扜V�d�:���[�h������8c�����]\�� );䈪T���(��k��8K"в��'�����ǀ&��Z��1��`O	H��c�!�u@��z��h��׊����"DL=z��ԙ�'� ,""�	:ހaK��<�F`2�'h4y�%I�74���P8H�Y��+�m�"�Pk�l ��A�;�OAA4�<߬Q�Y ��u�F�	|�����Hl ���%�_/z��@'�.Z����~���q�V�I��⟴�V�P�qUÿb���zԂ7�J�(�"l,�����?EVD���Q� �F��Xd�bcϧ%[�K��--pI�aH�e��]6�'m�����,5@M�&^�a�X��NP���)�R�.r���5����
���?��O�%��y�QN`��H��#u�����0bE@!�5D�x��Z5?L<{���~��8!Á'X�T��ű#F��D��:X�e�K7�\9f��>
�9	%�q�Y�n�~9X���ط V`��'/�O��uO+���Ñ�w��"�Z˦�Y�E� X�13se: ���d��%��	���17o��&�d�3`J\�����.L��a�H����x�6o;0,`��A.���2>�N�x�`��"���q�JO�B���wOx��@�q�&l�S�כAP��`"O�X������Z����N�\�=��"O�EcT��|Ld���a�.z���"O�����M�T�S%ρ�3����W"O\e�T�ٸ6���ЬAL�Bl�"OJY ��^,����͉h��r"O� ��`��J�"���C�KJ4jr �C"OR<�0��mfF���I,	p8�i%"O����3	��#��b[����"OR�J$Y�QW�	�<��i� "O�!Z5���3� ly5���%��%��"O�#5MO�]b�\�$�mC���%"O���4��5�T�D_� :��"O��ZU�� lF�QÊ��(dL:�"O
pu�̞u���s�E���ep�"O	��^��9f�ǏU��� "O�qD�I�a/���7A:�@�b�"O8����֯!�°��m��CR"O�� N4A2 kS�[/� Y(R"O� �eO�.���)��;���"O��+�-R����e��~�:!"O�Lh��L�T=� h�MC�8ɰRQ"O2��Ã
{�%	��Έ/g�T��"O��h\�[��jgMZ>d)�"Ox`�L�:�Nl24�@7}E��"O��k�aE�XNv-A��ʅ�.-��"Of�:�d�-o�H�0@S�V�Jp"OL(�D/���6���̃ �Iے"O6̃Ǯ�%SْmȣF��rh:G"O���'�!d,����=)���)a"O�)&�~d����+~�e��"OV�"��Bb^>d�)3
����"O�Ҁ]�H��䒗'�)�ܜ��"OnH��E%���+��E [��"O|9�ňپJ�d����3w<l���"Oܨxa�@�~ܸ��LU�'-P ��"O��.G(cڜ�3ClPk"�Ī�"OfL�����Y����K�o��
&"O���F��K>�YCJ3.ސSV"O��B�&ԟ|u��˅h�D�qS"O�p!�g����0�D{9N���"O�,b��2]���?0\)%"OJ�� �;\�\ ����\�ސ�r"O�sj�l�@@s����t�{F"O��!GI�r��yX���-��U��"Op�{�5+�x<��˟D�Zi��"OD��"OaI�X� X)ò���"O(\�1 �%��CF��+�<�)�"O��0T��VJ�{$��p�&"O	����t�xɣ�)B-

�:�"OezUr�R��F��$Ty�"Orh�wdS�Zu�=�t+O���6"O\|3�J��^֤��Ɍ-$�� �"O�qbЀY��*찤�Y�Jl&Y�P"OV��f�տ�01Z���sd��@"O�-q��!PԌ��V�E�Z �x"Or4�M��E�p 9d
 ?�I[�"O^���J�/x�M�������q"O���6E�<����Q>mҍ�"O$р�H���)Vē�I���v"O\$�!�ڇj�d�V������E"O��s6���g�d��*�R"O(`����.Dd0k�!�l���"O�S�̏�oƮ�v :Al�q�"O��#�A�x�)��	ݹjn����"O8�O �q�q�I�H\q�"O����g�p9�
�$zX8E�'����Q� *6���f�ҹ���d-D��s ?��l�g盪O�E�G)D� ��j+g��@cd"�8:�l����'D�� za��	k�I��`��YS�"O�PiReZ6��M�C��bb� �"O�4Qe��vY�$K�J�"O�l	���_p�f7�0s"O��s�O���d�{�O_;N�9 C�$!\O2)��Z4.H��K�G;p��D"O���J�I.*L*%�}��5��y"n�zj�y�� Z�nd��.
�y�ðl��x1�5wPasdŜ�y��	�(����O,�@�q�ѽ�y�]?U2>��5)��I�U��y"��I
,�cb.P�/��(˕Ɏ	�y��O�b<#��]�q�|�Bu���(O֣=�O�:ai���8�P<���.��),D�d*q�c�IZ 4ض�Y��6	r
�'x�dq�_�zr�IV�
��P�	�'���s$	��=��cU��R��'��=������Z�i��1R�!��'�@H6�J=��:ЌN�.C쥹�'����DD(Kxa�fON�-�Q��'�u����"t9>]q��®$����Op�=E���W�aa�d!
�(Nlܠ�J�8�y���@��:�O8z�
q���yR�,W0A�G']���ᇥƎ�yHR�x|��qv�i��i�[��yb`+e��E���X$g��atK��y�nvg0A�4k��//l�C$dF�y�I;:�v ���#�x����yB���Q4��DΚ�+��rf�
�y����J�]�b��Ӭ	��ܔ�yrE�r�R%��,���ӆF��y�����b�+��*�J� �W��y��Y�"�V��::��AS�MX��y���E
p��cޤ�5�Xk��B��I�����չW��T�!A���nB�I��x+*n�n��&��f��C�Ɏ*^BI�-I�^�PK�AS<qR�C�9L[�DH�&4{�8�
��O)'$�C�	/D9��N:|�
���C�# B�ɟ"���K���,���8�f��x�C�ɕ戕�Q�[�2��ుo�
&݆B䉸y�U[��i^�0�e�jM�C�I�U�h䚵��+8����.͵�@C��4��d-��N�|��s@�7��C�ID�*d�Ʉ�AĤ���
H5M̠C�Ɉ\'�%�f(5t-+�mDsƈC�ɛ6��@�r���i4�a�"l0�B�I�<b8q�cǛ��(��s�@-?�XB�I�XO���O����Z��ޡdgLB�	/�,�J��1	+P�m�_
������0A�%�2�)�:q:�5&�.D����	6[v����E8<�~Zfk:�Ox�PCf��tć7]�Ԕ���t�ִ�ȓ���	$�a��E���M<��I�+C:t�EpԢ�$�dхȓ"쪵������c��l�v�Exr�'BQ�wgK�6���A�{��!
�'�$�h0� c�mk�K��w��l��']�t��̑�@�a8'��$�Hyr�'�P{�)Q�s6^�C��P0'~�DY�'"����N(`�lHu��솬J�'O|�k�
�70X� 4k?hʕY�'�nD񷩊tD��K���}	�vO��*C�A��udH�
��a��"O�  �
/���'N=+�I�q"O���.�#r�`����M�J��"O�]��@�:AZ��$_#u���8"O��ԀV�g�*`�
Z����"O<dYv���d�Ë/]��u'"O�}�EL��(���Q%Q�k�z٪�"O(H�ӭ�~��s�܈)h�0�"O�ܐ�ב@|��G&��b�"O��b�#��<X仓,YD+z�Ѳ"O���2����T)����4��"O~y��F�=p��P',$���"O�����>E�X�暿R�	#"O��0D�m\�@p�N T�ޥ;�"O�*�,�Kn�m���G�.�*8�2"O� �<;�Ա���x��E�"O�]��쒛v�q�� ���"O
�ZÎ�W.J1ڕҟ4�ȋQ"O>��A�ʻ(�NI96N�N��L��"OT$ �j��2��#ߣ;��Dх"O�}!��#%�Q���'��r�"O��)��-��0!�$��y�"O�uhRj���%x�`E����"Ovh�Z�d��M�@����A�c"O>t�#�`�<��,J�]v
��"O����Wm�0��C+�1Bs�x �"O(EAՃ����A�Q'ݩ
����"O�E�m�)�J� GBm�P�"�"O0���txv��T�G"&0 �w�'�Q�и�F7 /v�+7H��?+����4D�l�u��-��qGɇ3�0I��=D�\yw�,�*�](eZd�0d�1LO��䉇�xd���ϗLD(	6�.D���GOG$ v�!IG�ΗW9ހ���+D�H�g�Ƽ+�=����p��`�g(D�Ty ԃ^�2�y�C�2$9d�{�'%�$(�O�I �iόcR ��G#H�XH�$"O�l�QHO�nq&�*�L��+�B@�2"O44C�n,��,:���� S"OƱ�i�2!i�p�!b��u�ݓ��H8���ҷ{�<`p�]��i��+D��P�B97��Ia4�[
��9����Vh<Qn	���%�4a��~����R�<��I��<T��		��YB�f�<A����.�X��o߇s�L���_�<yV.R�s��H�3� #P�@��o�<�Uc<1�J�g�U�+��U����Q�<���>S@@�C|��a(�HDy�<��$�9,�Ĝ9uHT0톅���@�<���%dM�5�ߨi9l}��WQ�'.a�& >K1���r�ѣE�֜r��׳�yBKʲ�� �"�R*��p�kS$�yK@�����N� w���AQ��y"�y�`�t��h{6�HVˁ>�M���sӶ�d�'E������5?���x���A>�١��3n~����KE*E�X(pG6D���e/�;G�l�U��o�FTH��8D���*�3q.R����7b9NQB��3D���ǧšp���t2�Yr�.D�8��o��©���7>�޹ۇ*+D�D{�Q!x�d.��"�^]�Հ,D���4�L0?hX ���0CR]�Q�)D����,��\iț,�:)A,'D����� C[4XNZ/z?�u�S�8D����
Cn�C�֠E���H�-5D�� � �q��C5�3�LW8G��m�"O��2vp���Đ�\�L�"O�(�7�ڳFm���p��$��aئ"O
Up��A�
�����
"t�r"O����m�oj�U��� W�d��"Or�S��G���}{��K��9"�"O���Q	�8Car���f�:l`b"OuȅJ��X��Q�S��%��q0P"OP��5�^��Rp�	tY�%"OL���Ǫy��59@뇛kr���"ON���|q�עb
ny�5"O(�,�v�tu��Ѓ d�h�"O��i�e�� ��e�8O�	�"O�A4��b�I�p��F��(��"O�,P�Pneba�#�G�-�"O�]�#Í&�D�q����Y�p"Ov����	�L�Ƌ��yctT�"O8M�K
"V]���Y�CLT<�S"O t�B��'\v��EKJ�����"O��xх^*�B���	Ŷ��)2�"Ox��D��/�p����U��4�2"O���C��7��p{�岈:"O��&ɟQb�"�ϛO�1R�"OƸkE��&�04�voZea�<�'"O�ԑʗsՌ�q�Q�/�ֽ��"O�I�cf_�X�2m#!���f0�5"O�5�7%N!p����߉30L �2"O�5kAJ�8
��lX��D�TJν;�"O�z!��$�@�Z"z.�� �"O��A�K�D}6�a���(�
�§"Orp�mH�S-��j�Z��ba"O6T�p�0d����
�]dr���"O��Pu��)?�8BgF�u ����"O�m�˂�<�����$¦��"O�ś� �XXf�[BMW[��X�6"O�@�qȯVb.<ZW���g��"O��@=M�X�*�n׵R]`k5"O�l"��5�ZR֬��Eo��S�"O:\@�.ܓ4{F�Q���5
�"O.|) �Z�yXHWK^z<�F"O"a�����;Z,IH��yjt���"O\�F �(P��4r3�T�\R΀��"Oh�c�˩4���B%$.LU��;�"O�} P̂�A#�����H�C=�t;"O2�+�@M�0��|;b@�tIL��"Of�cA�Z)��W��3$F�H2e"Ol�
��Ja��u+6��.cAjI�""Od,ij�)j艣��"b-��p"OP!*sŕ7\``M�r�&{#��c"Of�`��	R+�4ꑫH�I�-&"O���+-��!�vhЌ\��A�'�<�c�
ÛE��	���۶�+�'��dzD"� ��T`��K,e~@,:
�'p4��B�U3��0@��4Q���J	�'{
ٸum�%�Ԥ�A���D7��9�'(�!d.مr5�0+D�-Ϟ�c�'}��h�G�;Ds�T�AȪQ�!��'���ˡ(�^�L�c˕ΐ�X�'��u�S��1'f`ӂF��*�j�'�J!��#�ƹ�.>*�����'�N�Y����9gL��0$�)�&,��'�����l3-Y��$A��p�(�'X�S'��#p@h5g�*q���'��0�����:�\eXCI����hp��� ��X���9a�v��b()�j��d"O��0m��d��D�`�ݠp�n��%"O4���m��(��R�����C"O��`mF�e6ر�p�n��Y�"O.D C��e�~��U�'M�B�"O���i�+�&���I�!"O�d��Fϑ=���F"�9 FhY�f"Oz�a�k�2<=56�?B��T�&"O�����<wk8[7��)R�a#"O�I'ȋ�g�Z�a����>���"O\]�B�|s�8q�!K.���"O���椕�4�E�s���m5B���"O �0&X�n1XQB�7J0�7"OB]��$<>��UCT+�{*�0"�"On�0�jٛ2Gf=��)��P�f��"O�%�	�Mn�8�B�+@v��2"O�9��3x��=+��"A!ZE�2"O6="QN����`-^A��"O��{���4R�e��"�*W�D��"Ob�;�"Sv��`!�l��@0S"O4��p�Խ�鳔� B���"OVMa5������G�u�&�S"O���a�(��H� +ǬZ��{F"OHxmC�_�|8�#��7l���3"O�(�`E�D��MZaI�QV�q��"O�#w�R�+��p*�e� 4U�Y��"O��!���3n�)ʭK�1H�"OF]����E�^U��+2e��4�F"O��3⫊�,	�HT���x i��"O��Js!�*F�pEϋ�`���A�"O
��Go� t4�iJ���jHTd"OTAH�GX
v�`�/��f�$�Ѡ"Ǒ��<s<��ȕ�Ȼ8}�� �"O����X",�"	���*^H��y�"O�ay�H��:�d������ ��@"O�`��n��2lL��bp"O�(���[�c�P�c�S�5���"O�U�5L��4�na�	{��4�u"O���A�ڭ.�f�����\%�L!S"OX2��S�SN��1��	Ru�A"O8�K���W�4�� �#���`c"O~�Ɂ�̙y':��5J�L� ��"O�eR2�п����Q��iВuj$"O�yA�	?��@����u� <��"O�L�-�
����iV3;��}��"O
9t��^��	(��[�|����"Oh�R�\�p���B�*1�����"O�E�T-����f=۰"O8�B�&��[����{j̑r"O�@)��oF�b�/Ť.JUZ�"O�,z�,OTI��&,>Y��ɕ"O�Đ��Θ���%FL$�
��%"O.d�%.�<���c3�.��$"O�#�	")q	q���?&�ܹ'"O>,rӀ_�h����R�
�2T"O�s"�������3�N���"O�	���:��m��W�5�xՓ�"O�@W�$(�њ�˝k�B4`"O�5��)+@(����{T0�w"OP�C-� =�^��3�I%\N�;"O*=zĤ@�F@P����� RR1�u"O��cA��7|Tr�6���P5"O@��$
�|?��"#@3� ���"O����� BH�aO�?T���"O� ��s,��z�nA�ϔ��	X"O��z)F�9�H�Z��M��"Oi@q�
=��hP�"t��-��"Oā!��Nk�Qs� 4Z���3"O�aK��&@��P�҄/cz5��"OL���,�p��^6�4sw"O֘	�ϤX*=���;>6R,x"OR�����ʐ���L�B0��"O�!qv��oS�\�W�+P��$ʧ"O�� �"�"�����51�����"Or�CKأRL�ĺSlkƚ�(%"O��o�:%�x8��D3z��u v"O����H=v�襂C#���r"OLXQ�L�?#t4�sb�-x(��""Or���$��B�L9�U��"OF��0�G9}XV��O�u����"O�\��܌ʤ���  Gp�=�w"OX9��	>�B�C�#L@k�l�S"O2��1�B�\uR�*Q��NWd�"O�`P���5������	-0ڝ��"O�$;e+R�fkj��cU
m�xՊ!"O��JrG�ˮ�@�0
���"O�y�6�V�Q�A˟x�T!3%"O�B�@��]��jY�n���"O�$�%nI1���h�e�NA��"Ox83���y�(�E�}ֺ|�R"O�D�p�Ź*^�\��a3^
5�"O��J��ڴl�:���N��[z�iq@"Ol�{�"X A�]h���M�n8�"O�Ab䐟wc�Y����B��t� "O�8�Fb
�]>�E&G�l`�\ɴ"OTqIêJ������T�{Gz��"Of�1���-t����FB�b*\z"O�	�`�^�D��U@�!� -�)�c"O�e�G�+/�"���J0e@l��"O8��u�R@��cꏚK��}�"Od�� nE3��s��¶	)RqQt"O��2��͙B�\�B�%�m@"O�<1�!ϊe�lHP��4��"O��P0���10�]��FJcה�(�"O6�Q禌$J
2P�Fé"��ee"O�mʰ���dT$P�"h8-CL�y"Oڕ�%�*x��M���!yJlY�&"O|(�f� �3b|s���D�~�)�"O����C��W��)8�"��8�"O��[�E�ELx��@v*$I#"OVā2�΅@rְp�E$k�D�ˁ"O�=�7�
P�3�]%�0�á"O
��@��d�^��A/�!Jq��Cv*O��@�M�.J<a2��`�����':L�(6��w暐;҉�-g��HR�'��x��V���#�F�W�^��'J���ۺ{b@��L��hD���'�"]k�-�|ȸ� m\�&����'<�X@&�]���¦��nwyj
�'� $K3H�B��P(W팻5,@�C�'&�p9�j$>g�(���0L��C�'��s����Q�C�K�O���	�'�`e#�I�)X*<��ZY`
�',
�yց����q3ܐ(�
�'p�ܒ�Z�0��8Ԋ:�*0��'�x�sA �?1����`����:D�h��9U���qD
$�pd8D�0���jK�
�M(4�$��+7D�� ֈ�b�:^s����D�F�)��"O�xk$I2%�>�S�E�1�Ρ�"O"�� ���P�D��`��y"O�Z���).K@P�"�+��{�"OL1����v=v(��8��T{"Or�Jrl�ǜ V�᳔"O� ��I�0X���V�R-2�'m1OL��֏ܲ�~l����W�i� "O��bd�!�����\A�~�4"O<i��nO�"#,�r���-�miC"O�L ��C�
0�S�b̶W	8�"Ob��e��}��eєO˃b��q�"OLQ�Ϝ9Z <jp�ȗT&P7"Ol�"N�I����Ŏ�,f"H=B�"O�aQ�����(E�¼y6@�6"O��D�L�;�f� i[5?�$i�"O�Q�ԫУ7kd�� "�w��d"Oɚ0�փَH[���2r��5�"OhP�ӑ|.rA��O�(,L�6"O����M=�(M�%IH�(���1T"Oi�!刕>l��+��DKd"O,E�ER��%qTgU�i���"OJ�)�.V�?TU��E.��1;�"OT)���  x1D��Y��Z�"OV�Qc��������!y(�0"O<���$i�4*�`����"O�Q
pLׯ.�<="�F�:S�H�'"OP��G��	C$ձ��\�=M@��"O�@�$KM8u��A!�l�O4��5"O~�:��V�&����Ꞵ^��7"O, �3�ь#��q���N PD��"O�%�q�R�|�HJ�`�����"O���1�

`����P�����"O�9�)��0m0) ���u�!0�"O�H
1��"(  P��>��ZQ"O�Ԁ���~�p��a�� s-�,�3"Oz)��&,gȥ����.\"
i��"O�58�A�}�Lc�A��sRB�	(i�P��¡�&h|��1"	P
�zB��%s�J���D>.N���w	L�Pq�B�B���u���$�밨�'4��B�36�����$���!����B䉋 ��M���*=B*Ya^>�(8�"O��ca��=:�xY�h�3$(Y�R"O�h�3��`"����ڂb��pk�"O�APbR�(�ɴ�}�d�� "OJ�Pf�8b�.U!ӏA2�0P"e"O����{9��	P�ҿ����"O�I��e��A�W)"���"O� C6��)F%�<Ґm�� �}X�"O�*W�$7l��Ӎ/�"	"O�@���o-s̜3h$ƈ"O �#�ؒ{��@�Ũ��Ԡ""O��pu��@U�Ԋ&�4P]BW"O`#BҞ1�|�ɓd�#�>ei�"Ov�6EN;w�|�9�³h���Jv"O� �,y&,��	61�����`�<р [�� �[R�.6?�ɂ��s�<�$��$UrTy#P0m��1d
EI�<�We�x!��L"w�B�Pa�F�<� 䀎�ʡ`!�_bnz���Lj�<����5n �	1%>Ŕ�2�j��<�a���1G�o�Vēqf�F�<i��
%���a�ʐ;%��K���F�<� �Q�6c¾}��MR&�$�i"O����þY<�`��۩���"O����
����UAz	r"O��wE|�`�`TMH�?#j��p"O�P2Eq�P��櫃+>���"O�	�C��E&�L�W�B!^q#W"OqY֢#턘����R�z�"Ol�sv"p���((�5�lږ"Ö�e�6=�"u����),����"O޹i�����F��Fv2��"OJ)Y�&ъ:�m��?Sk*���"OPɳ7# ��X�j�&|��T"OL8�W�+~f �ns�
iX�"OjY�K5i����o�p�$U��"Oҭ�#�� $��!�i��S�l�Q"O䨫2_�|�ji���M�
b\�q"O���eiͲ��i�B��xF�ٚ"OH��(�R���X��ËT2�E��"O3��0���+�EOv'�ܛ�"O~xee�9=ҽr�	.ց��"O��*B�K,|���rA�8��q0"O�`�&�4f����E��\�4"O��÷���!�� E� V<4C�"OP`�Q���"���`�&��O�6��"O"����-2W�Q���9=�漩&"Ob����R�U�r�h1f(���"O�p؃�F�i��er�&�y$��"O�}��#T��J$&��y�F"O�E��Ó{�֨���V|Z8ks"O~�IҬ����7�
5��  �"OTh�%�O�Hڤ\)��\:{F�;3"O���<�h!�Y�S������"D�@�@E��.�8�,H��ĥ D� ��OUI��XQD��/C�̴Q�?D��l��F��&C˛2?��U2D���l[E��9����J*�8�5�"D�� E�3D�H1��U.�Є)Si!D�Б3L�,
q�ҭRb��"v�;D�i���=FG���Q�Y`�E�p�9D��0�ӃX?��hB�":I�4Sc"2D��;��N/R2$q㨌-NԦH���/D� 2���f�`�d�J>DUr$"�e8D��h��Ҡnt�"c,U8h��An0D��A�HVN�x ��.�l�*��/D���A	��i�I:�ꏰ*8��0E#D�P��L�	G㰔Ӧ��Jt&�A�� D��x ��,a��{�F��a�����$#D��+d�P�e�tP�eǗ�%
ܑ���"D���R�E���K���5	e�A�En!D���eC��YX.A
��}UrE���3D��q�+�=-xhp����h�Y�`�2D��HCE��|N$��k�Lƶ�)�+1D���W�K�y�&!H�4�`l��H/D�l�$��5�H�s�䅡N�*�P­7D� ���.n��p�Q�O�<*�(ah#D�X�G%��~_(`w*�3x�Щj (#D��@��V�t�g�������6D��{W��)��H�,�?r��$�T�&D����;Q ����?1 p���!D��
�gӼz��E���\`A� D�\�T���	>+w\��g
�0�B�	L�FL��>
��
T��7(C�	,9��=S�!އ <��A�tfB䉫#2  E�ۏ�h�@䇔p�dB�)� �IY n��bd�l���/<�I�"OnQ�iV ?m&�Ѱh�.44�*�"O���w��Z�Z���[�0^ʀ"O�p"
3�n�Q�'[�_df�
C"O�Cp`K��"S��'e�ijt"Ot�f�Ź.�0T�]"�0��B���y�mIP�����HF�z�JQs2D�$�y���'?��D�W��!@P�2BÌ�yb! 0CP$ذOC2fÖ��a�	1�y�n�gP hC�^Z2���pd��y�šI������J�I�Z�k%�����?��'/�1���L̩�Co߸>�D��'�<�HAHA�B]�$��
ʯ2�Н��'���2�B]���3��|b�a
�'������R��J5����U�<�Sj�_�� PD��
�c2�N�<���}���)�&��)D%s�a�^�<1	�옊F��>9`2�R��Y�<��EgN�y� �H6��� �W�<��:='�i���'\�=�m�N�<Te$4H^�s7��="�sRMH�<at��V����$e�8r�B1S��o�<� �5�~�đ�@�4�0�GA�<)�a_>��v��TᐉQ@�<�t���e1��+��#H�*X�%@z�<A��Fz��dL�9���#D�v�<W�ʀY~`��?W���Hu�<q2ѕc��	`f�=6p���D�W�<a�8'�]2f Y6@���{���M�<�C,I
3����߻&߆p+GK�F�<I��/������J�Z��4����f�<q���1�x��`�Y�'ӆ��f(Zh�<ɓ�D��ԫ�(_�[��p�h�<ae��#.B8�%Y1TJ~�jS�Eg�<��*�s���`O�Q�8��[c�<��5oٶAs�rXl� [^�<�WDR8K��Q��!����(�X�<��(Κ���pi�B��wl�<��Z=4�Ȣ��]�[����Ul�<�@g+�D�S�j�F�\��t��o�<i0 ,s�BQ�CK��#����fXh�<��E�'u�ȰFm<���Kբ^b�<9h�|z�$�@�١H�1sgb�<q4)kײTFE����ِ� �y�<�D���*wĚp�^kv�<�mƌ1VԬj�ԡ���@� Fg�<a1�V�
����:�p��5śY�<a���@����@����N�<iv�\�+�|��]�|3��03�@�<1JZ!rI�	� kr�!Fl_{�<��
Y5,�T������V�8���u�<a��G�?ql������~v0��g�Do�<ѲeU�G��D����x|��[k�<I��a����po؝e��)�|�<�!�ݒ.�D���Zu�� ao�<1�i �j2v)�B�}�Pi@ǃ�U�<!1��!h
��`�A9��	�@Xh�<�3��<��E	r`�tR���c�O�<�G�!:P�T]�H����H�<p%��~�h\���T3x-��ٴo^�<y�K5~f�U��`����Հo�<��	g
T ��c�(df��0©�U�<񦨟m�<�����!?�ȑh�HJR�<�o�>s�8����kΎ�ӆLX�<� �ñ���q� �1�O��Y�=ra"O�I��f�O�D�9!�ȸA�f	�"O���-6mc�)��\7nϰl�e"O�P�R��F��6�ڣ{�*m3f"O���7g��Ԭ����e�
�'�XJ塐0�8Av* ��=��'8�1%��Wn8�y�
�'NL���'�T)�t#ؚRވ�(��M��'@��d0UV��Ѧ��_^p
�'a�4ab�O�ly�@Ȧ(ȭ�Va�ȓ[N��$^�q�F%h %L��=�ȓ&8���6�_�rH�0���!H��ن�O��8�H�(�}��KM(LY�ȓ�~� �J��?��LH��ԿH�@L��J�l�w.�:w{x�	W�
Jv(�ȓ(!��k4(ˇt,��	��@�&L��A䐴��-�3oJ
����>!d��fg^\��g�6*|�ᢥ�_�61��ȓ)�Z#�H�ef��b�.�<#�ɇȓ@�>���S@�
pB�m�����	Z�'����UaP�������=%�l	*�'�jx�_��q���B�n��)�+[G�<A��(��� �t*�W��F�<��9+NX�c���{��!%�<��J�e����bj]�I�����x�<q&����p�ܐo*��m�<��F"p�^�t�D�c�̨��l�<��*Plh	��q&9P�-�g�<���K YgT쓲�ܒ�*�m\]�<�@�W��B��(8ȕ���W�<��,Ӷih���O�t��M3%�W�<���H�=AV�2Gl��9�P`Zю�Q�<!����T=��Ƌ$��="CD\Q�<	V͉vL��&���\�V�a
�A�<A��::4|4��A�842�Ui�<�g��}kR塦I�0����`�N�<����b��\�q��F�����s�<�j��a��,��cA�buJ��@��m�<yvf��o� i6A���Y� ��i�<CeWGl�u�M8n񢠡qg�<Id�#Ab]��ˇ�`�q!���yj%��p	q��*-0|h����y��;yv	r�J�:!16dゃ��y� ~}:Lx�(
�C��\�"���y��T�gM�8���'P���Z��D�yr� >/�� ۡ��E)��ӕ�Y��yr/��d��1�ʓ+.���@e�\(�y���%<Є��ߤO�z!)E��9�y�DU'kn�t�ͬG7�
U�S+�y"�_�Ka�ax&��U�����'C�y�b+L�&�Y���>F_p8B��y�iH���,XT�ĸ<�fm0��y2�I;Z��"��5��Y
B���yRY>t�.�óGQ:3�@u��=�yR�-<�K��$���AHJ��yRd�����5�� n�R�'��y�a��OFT�'Ό�=�Z4R�ک�y��6@Q`�S�b��9����G-_��y��[!I\2�A���)ˈmA���y��G=�\0�É��J`��A���y��>X���"a��yz��!�y���p�D���	�f'�IRB����y"�V��U���M�^m�ˑ�`/D�x��*�WAt�r�T�l��/=D�� ��R֬X�F��|jC��-g�,٣�*O<��S�.|�ȤI��F�L�@���'�$�Gg�:C�jQҨJ-	f�s�'�8t
dk�[ې���@J��C�'�Z$R�� ���Zt�U1~�����'jl��U��� ��oحr6޴�'ŘXA�ǉ�A���H��c06p�'�Q�
&��i	u�A�HD��ȓ:����4�����5���Y�A�H�ȓdӰ}#Q�l����7�^�r�⍄�����Ph!��aFZЇȓJ�4�s��ӃD�T���W�R�Q�ȓj9���qcХpDL�a��'�ؙ��Y�n��Ro��κt/ʧsRY��Q�n��ՅՍqFL�е��PS��ȓ.�p� @D�L���+�"ǣc����ȓ
wp Ib�B2>Ɍ�� ㈟=���ȓ3hqb4*�n=<�d��a����-a�+B�ި[�P� �L��/�`��|�XT���������g��(dY�ȓ4$ɺ���T��u�Ξ+Z���r|�X�@�L�z��b���wv���ȓ_��iZ2I�%ME܅�F(X�[
Rч�#�b�
S �_��R��
�$���ȓ@��;���"*F�9� V- t �ȓ|1P��uD@��%�7�^\�ȓCKL�H�H	J@.�"k��rE��5pZ쫑!L�4�pX3W� T����ȓSl�&cV-�V�����;3Є!�ȓ�`a�d�3
�=IրZy�X���>��q���&v�Z�3&\�d�ȓP�(�!ѣ�46ތ0R�n�q ��
�l���`�M��uh!�WH���_pbY�/�e�V 
Ѯ�5�:�'X�<b��H1V~&,����a�p�
�'����Aa���Fe�3�2W0�|	
�'ˎ 9l�+��-��1Rp�1	�'S�m�/XF�@y&��w@�	�'hR�!�+�� �u/��t�(L�	�'�B9�� V��)j�b�&W��A	�'�xU(����2T"�jǩK��i

�'T|C�jG�o�أ慙DX��h�'��j&/���(+�H�5�f�q
�'�̥���ӡ=��9��4Q��3	�'�a���OH��h���+����'FYbB�5�x�#LʵW�x�'
�B$�dH�p�n�|S����'i\r�3<���	�yp,D��'�V�)t�$?�dԁ�kI*v#��!�'����aT9Ӛ���,�a�`l�	�'� Y�"�͈x�8 �6���^��A�'g� �K]�:%`ٶ���PI����'p��!%Q Yިҡ ���'C���hK3&�]jr�Q� ����
�'��b�7Y�$�c�C(2�L��"OP5���@z0U;�gȃ*�(��"O�)X�!�(��Q�p&��p���8�"Ord#�J�#.�*�a��8:MyB"O~`)BaO�1�����1z�P�"O`)y����QG�&�N��!"O>�9#
�H>5�B�q��D�W"O�����6�T���Z�8�#"O���P��x&V�����F�^}�v"O �ߩ[~���l)@�ܴ��"O� �IB�I�v)� L]��L���"OrM��͌�pY�pI�Lk�|�""O���H+]�H�Ňɮg�c4"OF�KK0�z���E�!q��"OX=W	^�k̎q{��XP��H�"Oh�0��.#v�� #5l:��'"Od��gJ_�@���a�>U2��"Oz�(��	j]��#�{ ^	�%"O�l�$�E�d�5nK�A��Ȇ"O<k��0?��+��BD@��"OT�ZZ�|�K�6,��ң"O0�H�A��	��e/֏�ٷ"O��!��.n�PL��i�b���"O�|���L4%	̝K��I�}&D�"Ox�b�%N:wt�!�a�+P���"O�̒�N�פT�pjO�*��i�"O��T�͌7.`pv��$�G"O¬Q#͘�b�U;�N<t��qr"O �� F�
k9��)��ľ\X]��"Ov��ǅ��F0���h�;B�r�"O�Ӈ�ȭl�zaP�f�9��QCa"OR�����E��]����c�`M�!"O�֛}l��5�ĸ!�"%��"OV����Y�FL�C��޹zН�'"O � !֥�8M� �ٜJs�%�"O!㢎	�`t�d�46���0g"O����<6Β����F�Ó�7D��p���!!�f�U(��U��	ze+6D��R�� ����Ńp�HM� �2D��II��/���rC/)8n���0D�\25J+5���%E� �D(�6�.D�$���t��D��H^�Y^��y#+D��i@�v�*�x���G���z�*D�X��R��,�ŅۂuN~��(D���u�\�3�^UhF�[;
$
�C��3D���ᢆ���iSR�Z�Cĸ���a0D����&�3$f�i׮�>;�Z��c-D���`C�[ ����'�~*�Mp��)D� #ĩ>#
|�䔏,�����!D�l�%#F�S�����a��5P����N2D��!(�-	�f���$��|�2 ���"D�4�Eoƺ�n0�d�� ��ӴH D�� �6*�B�H�2�A`��9D�9bǗ�"��fɫ46��L+D�<z5���X�b��LG�"^2�TJ+D�P�qֵH"�Q�#��&!��=D�p��+��,���٣���x	 1� �;D�,��
�M)�-��5[[ �s�7D��$Lʹ�"Y����7L��{AA5D��Bf�%c �sҌ2 �:#�6D��� �\���0��ђ|\��� � D�dC�$Dx9qv�>P�$+5O=D�\��
?�L�He�m(x��m-D��*�
��tu&X�wAŨ&�xQ�-D�<)�ޠ#Gf4x2��-Z�( e*D����R�{tx����U�h,چ,'D��h��Q��`Xs��:i���a&D�xQG�5K��I�	�Y	FeJ5�%D���T���Q��͉'�1��/D���ێ�T=��
�(���)�� D�,�e��3{��g
J4/|U*�3D�Ȩc� n�t�hQIH�o�TE2'I<D�c��V5/>�QD��~>0V(D��+���9���C���<[`,�0��'D�� ,
�	ҋG���]�[.��"O�<
�Ir-�8���2}-�a�"O�3����u?ڵ;p-�)�)�P"O��1��+u�L����l}���G"O��q�$� 4���ǇL`d{#"O��v�����YQIMG<b�Y"O�	#P�}i,i�I� ;�4�"OB�X��mA�� !BY�`J~�)�"O-I�,�?.���f
R:�P"O>�i���,n����Ԅ4N�(��"O6��3�Ӄ|�DH����{Ӡ��b"Oz�CᘽS�������`� "O:%�Q�ܜj"z亡�_/aܞL3g"O�-���*rn%�@IN&Agv�2"OYa�V�A���BuBЯP��Y�"OF)vFL�{+��f�� !���{�"O�e@�S�tQSJ���h"O��q6�E�Yr��Ɍp��D�"O�|ȅh�T�(2�&�����"O$�@�� �$m(��57o��2"O��17*�	�j��&ˌ'`���D"O��t���1��lH�@��M!�"O4��Mۖ'��%�Iɳv��&"O$Ij�f�)A���AS������"O����ݲJ~�VA�c���#�"O�J3oE Knl�U� -����"Ob9��n�a�x�c���_u%�v"O�Y�q,G�{d��F��|.��"OBp(��F7K�́�f�8i���Ȅ"O����m@CJ4Q`��*�q�"O@���`]�AuJ����Ⱥ���0"O�J���&�2}�V�����qt"O40 ��P�"P��)!���4���%"O�<�s��D���񌛃>���s"O�9R���Ҕ2`E߸R)��x�"OPc�,C?c!��8���!j�w"OpP{*̷Y������B�[U���q"O&����uQ��)3o9����"O1��LБ�X8�u�ڒR=�i�"OR8��!�	`��o��_ ��P"Ot���f_�,���`�طP��ܚ�"O�e��Y\L��
C��]b�"O���&Nڎag�qc�nH@9Q�"Ozu�2$ʱ_U@P���@`����"O"9A-Y�oV�y�f�$5�]�W"O�� ��#W�L�V/�B�&"O>��OC��t��Db�D�%#e"O:��F�0��Ih���#{$�"O&D35��9,H1�,Vj��5"O�!���n�PX��{P$�S"O �*'�dH��f�{J0B�"O`UIckE.`�R �DH�&�=9�"O�+�JE�zc֬
�E�!1��"O8��6�u�PSeX���@�"O�(3�r��3�dΪD�ى�"O"Ex�)!A����LR/9-"��"O�!�F�'<��eM��1&��d"O�a"B�
L�Н���
$-�6�4"O��IS!n�v,�)ת�D E"O��aBV�7����զڕ�R"OP�`�غZ��(���.���!�"O\��kѐ#��8K'���Vm	�"On� ����iyGn�fn��`"O��z��]�	�FQ�V��ljF)U"O� $��V�{`P(�ǻ~�C�"Ojx��˜Z|��F	�(����"O�����!Wg
m�%h�2�@��&"O�9�E��Y���6F�K�,��0"O�%�ØaYb zPg�X��mY"O�S	���.�8�&�#!����5"O����*sA�$*���zVd��"OP����t1��P�c�69�z��6"O8u����
׸\2�C2_��%��"O:�0���;A�|��O1 �I��"Oڬ�Չ^3A�đ!6(Ճk�@�z#"O�!q�B��
�.��2-��<hH�"OB	��J���29�H?r�(��"O�-$��yK��b��=��d{��'�ў"~
_�Wj
`��`[�%��U ��ͫ�yb �u�6o�)ph���$"�0�!�K�q��!U��,}�~������!���.�f���K"&��x`a��+!���5�����	�I�*��ek�;!��	���2En�O7\��2C�!�L��9��mݢk j���+͏/�!�6]��!vOa&�Y���!�$	wI؈�ǟZ|�x2��K5H�!��k�41CVF�jh2������e�!��=j�6��0FX�%87�&0!�$��<,<����:nH��H�)�!��,/�* {7��fH��r�ؒ�!���'3pB���޶{X
E¤��F\!��Z�0�p�=�`����&�!�DZ�tn&�8��FN*X�kA�;v�!�ċ�R{��sL�=G#���f��J!�d�>��Z���%"���AO�T-!��ݞI62PpbaM�a�����G-$!򄉀J���{�V�o��D!t���:!�DH��d�`TJ�1jl>}@AL�/v�!򤒁V���[WlJ���mY0���B�!�Z�)t�2�$�A�dDL�<�!�D�;�P���d̳8W$)@���w�!�D��j�h����R�_;���,K�!�D
;�*�r��M�XhDM�Y�!�䋼&�8��g??`�3�^�>�!�D׼l5�����t�xɊ��K�0�!��ڣ6��H�$�L�@�u2#�a�!��-��I�MǷ������<*�!�$ϟz76��T��!��jeb=�!�dL�`�@�b�Z��G�d�!�d1�>�Hԍ���
�Z`���,�!�$�� �Šŭ�2���3R` �!�D� Ô$��]
fz
��l�w[!�D�Xf�H�F�)	j��@7��!.\!�d��ReظXĆ%lS
���C<HN!�$Y?&�\s�	,r?t�tmѸ?!�d�e�~!��P%$SWl�<b0!�Ā VV} �/��mt1l��l!�dS�A�X�����Xm(�'Kͩr�!�H1OX�I�&1\�� �i��!��\<�T�q�Ct�� �H%�!�A�� �"��U"��29[r!��A-���"�X1��X���<p!���6ʈm�d�^�"'ȸ��.L	d!�D�4d�R,��À0!�xQJ4(�mH!��H��5)6�D 9�'�4}ܩ�	�'Fx�`�)A��@c')��Y҄��	�' ��A�?jX,h$ֆW�B��� l蹳oɼKm�D�����Л2"O���3�E�~u̡�gD(�����"O�Z���)+�c㟅/� �I"O�$�B'̮7���6BQ �^�b"O�c���6�
L����k�d@'"O�}���D/G�ք"��*4� ���"O��r���V��X�ԍK#�{�"O~4b�/ 5�Rc�&�%�"O�I�VM��V΀�BE�T<�1�"O�Y�KH+6��@��3x���9�"ONi$�������z��љ�"O���!��U��!����^mD�K@"O�86�ʢ7{�pCDN�Di�L!"O
	��R��`�d��˷iC��y�_�N%�ZgW1V�^���S�y��U��8�:� H1a�����	<�y�j�:NN��HZ�ݲu����yBL]2H@��QŊ�t�ť[��y��
_}h|c��E1y��EZ$�>�yr���c�<ث��4j��L[d���y�a��$'@L��\$fS|p�j ��y�Ǔ!oV0DR�n~!����1�y��ߋL_�� c�.5�h�iҮZ��y�R(,V�1KR&R/*1�p�q�I��y�j�u��P1g&G&&ObDaт�?�yr��S���bn׬R4B�8d����y��(~$Y�揶5�L���B�yB-�,*W��8aL*0-�$�ׁ�6�y��_� ��(��Y��dpǯۉ�y2nN�kJP(����H�����y��u��X���R�<��x���?�y"nXʈ��jQ3��	�S��y��X�1kd��a�Sp�'g^��yb䅸H�dIE"���qJ��yraL'?,@ҁ.��H<��1�P��y�Y$t�bك���EØ��a
�
�y2B����Г�֞��yaO�y��|wνA�Ƒ ��b�&+�y�K_TJa�b�Ε��@�.$�y2��>q@ԁ#[�}�R����yr)8z6�k�E������d/ƅ�y�'D�u�z=0⃖ 6�AjT���y� X�BGZ�bR@��f\x����[��y�h�:S\�`fA�`�l�+2����y"kǧ$������5d� ���yb�G6T��x��Q�UǘD�cM�7�y��
�a(�*�)_��P����y�ۃmP�9��*@?P�t5c�e��y��_ �D�4��48�.d
`�y�ՏW�J�r���3���gl1�y�aIi�A��m�'{|�{,�.�y2A�cF�p+b!�!&�Љ��A:�y¦J�"��hIU%4@ʈ���!�1�y�5�F�`fn�	L��3����y�$nq+`��7�ڙ	wi���y"��.��0E �"@�t��C�yB%�"�V���Y�0h�Û+�y�h�tz`�	��!挅����yrʓ�<Cl�.�-�nN�N�D���'>V-�KL9�-C���$��q��'��P�,��"�j����S<f�.�J�'R�@ߞ'd�ɂB<a� �2�'��$��.+5"��Q���R(� ��'�di��Hܼ�j�#}�L���� ��ڤN.]u�Mp�	���Iq&"O�E�@@-�Se?�Rq�"O�4�סZ�N�\-:,�M�y`q"O�d�A�'k<12	�
J)I�"O�0Hj�'1d�-X�"O<�k�ȏ�K�� ck[cb:@Z�"O�m2$��-!����+��8m��B�"O�,@�MTp�!��ሂL3�xr�"O^��SlM�2F
E`��\�
����q"O܅�`�)<J�Qp��/?���3�"O� ��p����XwV`�1"O���nOj(CE�c*$�@v"O��0c���`��r U�4|^�k"O�-j�%�1�D��B�h>��jb"OD�b�C�ny�i��h�i1�a��"OH�H���@c~ـ'-�*��$"O�`Z�����u�L�T ��%"O����	͈��ǭ!����"OJ�:�Ä�:I~8�t�TK��Qd"O�J&�!|�2pRT��3V 0b"O\��S�	^2����UUFZRR"O��i%�J�-�y�Oٿ\0�uRf"Of���)��,�«ֶn.�9�"O is����/B�sA��j�5h�"O��)������A���O�"O��7�F	"4K'�&:���z�"Ox��H?X�Ȝ�G���y`L�16"OQ���O�/ʒ��.^&��C4"O�J���?\��҂�*L2
}Jg"O@cf��C�ɋ��Bh�X�"O��GJS?P�v��j�b��љw"O*�'�8?؞ѱ!oVQ��P"O�Q �$L$IK���/`��BU�,�!򤏝K�~\2�B*�J��j�(�!��$�\�aP��DT:D)��l�!���>(�C/á;�\� ��o!�������$��+t�A���H�o!�
���S(�l�����:��DI���e���<W�!�ψ��yB�E���c6/!Z`��y"�2	n�eЧ�)��A"�_-�y�(�<8t�y#GF\R����1#ڎ�yҥ؀Q={W�,N��q����y�3U��3K@�?�l����y�[1g�dڗ.�:��=����y���:c+�h�d��k|0@'ň�y2�B�<3\5�2f	Q�x�Iq�<�%IƹF4T���E�ܽ��K�w�<��H¢�^���p������w�<����,�x�a�-�}�B�K�O�|�<Y�C�OHxx����V8
 	�v�<���M�8���a��}����g�<��"̚!ԝ�cL�Y��(բ�b�<��H� .��Q6(';�a �.�_�<)e�[&{=b]��ć�xP}z�F�_�<���%��P�%dαu2�E�X�<�Ti$e���2����a��ubA�R�<��m@�{�� z�,G�7����RN�<	A$	�3~$C���e$h�Q2_�<Q%B?������r�li��Y�<I!)^�w��}Paf_
o��)�`�<ᡯą<g ��6��\�4�`*^c�<����5���h�ɗj���Q^�<y�z��9����@��ѻ��C�<� <!��(3�e �a�B{W"O��Ҁ$�M�<Q�C�]�t:NxXv"OT
v�I�YG�E�U��-��A"Ox�qb�o���FgVh��q"O
�x�kV;�m�e?<�B�&"OD�+��Z���b'�ӿ(T֐!4"Oh�۰��!YT�qWA�0V�R�)�"O��Y�!�j`C�O�z�%�r"O �2�]��Y���L���:"O�� S@�w���Bo�l10���"O��Q� d1�L����I� ��"O����L�
r�5؅�B���l�"O����̊TG={c��1|�X�C"ORt9ĂջV�<�����3 {��1�"O�<C'Ά�v٘y�B�*#�<��
O�7-�6�r�Â��$a+t��J�!�d��3���k�a̾m�rL���ջq�ab�O�	�4�A6v��Ӆ��-�,��"O��KC��[����%�G�'��I����3.�L�T�A!_H�l��Xt��B䉭v��	���ף=�عգ�b�Ģ<��T>E����'6x(�`*�!'�P��)�OH�E�f��s/��ظ���I�LD�9Zd�>����<F��'���u�E�T����p͍�?�|�"��B妁F��2	�ؙ��pH�-���V5��ā9���&�ē��'vͣ2���
$��j{��dGu�*@�?%>�KN>��zn,�q���n���a��t���=ѷɍ�_\�q���0h�������f?�۴���g�,����OG��賅�P�� p�cK&L��-��'�f��1g�+L��$z�	=Ib Z���'��>���2	�h�Hи"�����;B��B䉈j��H�#aY�g������9rm�B�	i���shK�x՜0��[4{0C�/[o�`�c��p#B����B�/%�<�g��-7z�1t�Qm�B�	C����G�+N������.H�B�	 Wl�%s������蘒U4���0?ل��;d� ��d���g/<�WB�s�<�"�X(Pb�)���C�i��D�P�H�<�Ƣ�:J�2��[#.�"iP��SN�<!����E���s-b^`w�]L�<Q"	G9?�nd�Sn��ǧ@K�<!�Tq����*�_�*�KU�S�<Y$�.���7gY�*��b�O�<�uH*aC�A�=W��(��-t�<�Df8����qG:q7.M��Yi�<QD�s�,k�jO�L���$m�<�vd�'��(�F�K�|�Y���e�<�֍�c�-�N�E�l�)5�V^�<���G1
upA'V�M->4z� �`�<9��ֲxz	�#��k���ykXQ�<	 ���0Ը��!u�x9$�NH�<����*zP��N�*�\��%�D��E{҄N qj�����5.Ԉ1�	���yBc��f��	p�bAS���1��%���(�S�O��!ꦢ��T�T2�k�% j���'
 �7	��dF<��$d��b=��sJ<��W��@1DXFJf�7�ݔ8�@X��k��:%癶u�,� �+�|�����i��L*w*��#1���H�E$��ȓHQP	K�FCP��գ�==���IFy"A�5辁IW����.8i3����2�S�O鮼�S�$tb�A��H@H5��EQc�']?i{�$��<���H�2�"��"+D�� ��jM6�~�xBM ���W�x��)�� �����!R�x�.�� J,�DC�W.�Q gΔ�H�ň�͇�M�a���X�������H�L�&d��O����杠lfH$��*O�2|.D�O$Dzb��(���A���4�{�׉q�!�DV�� �S�ȥa��ٙ#.��L!���`�-��I].,�͟�L��b��6�S�4ǋ=K$����G6_�بaJ����>�J���Џ�+>��Ӗ!�"�f`��JEO~�:O��)��<���;��-#A��� �:�#��jX���=!��ZȪָ�N�	�cA�8����O��M�
�x3���lķ[r�P�i��`�I�����!�'��S�ahW8��(G Ɖx<�P��H���87mٔ���)�Ɇ�]l��'�|�?y���B4sʍ*�E�:@�����ͩ!�>X9|]�c�R��p�W �6)n�ӂ�)���b��0+I, �����8eޤ��$ȸ��Wv|a��Թt�hj4+кu P�<�ߓ=k��ۢ���p�F��Щ�.2���>��'V�dq���O,��N<�@���^��d���I�t�!��K4*]�
C ��x�����M�铒��3���lc�����&fv^��$N&��9��6D��j�Zc�)*UŞ*��k��O�㟨���?�sA���t���<<QPǂ$D����%֭FW��@ϖ�
��5�&��O"�����S,�:4��X>�tj2I�.Pd��ȓ&�v,
���##(%zc�)lo��'�`���	�0��A�����H)����0�c�XD{�7O��u����/�RՊ�e�	m�֌�ȓi����-As�l��Ř��B���OM��O�-Gz�Oޔ���J��0X\m��Bh����+�I�a��D��AZ,���;����ɣ`X1O��G��O�#�퓰�,SVF�T.�\��"O���ֈx��TuNB�&�T:ѽi�I`X��JF� ��V�2��U�4�:�!� %����Ms`V>]أ��JՒ0R�铱n�"�z��$D�hZ'�?^T�6c'5����H-�h{�b�E�yG���d� ti�3���R�<�+��Uf�y��/�x�u; ��S�<Is��P�$�`��H��#�`�y�<!v�L�Z�V��$ӫV̠ي��Cq�<V%�_���16jSV��ܳs�Je�<)���)L��I e��+dʗX�<ɲ/��@2�����݀1i�X�<A*P�R��ѩV��?WJd	aZV���'�����v�� ~���C�i,�y"�#E϶8I��H6w���$iJ��yRj�Hx��p�D��"$��y"m/�t����7]L$)�D۟��	B���Or����ކa���f��\��	�'1��Ӌ��G���0FZ�
����';�5�'�ھh�$�q���#��ӓ��'�*�ʲ��[��b�T�U�Lc�OR����Rt:�!W�#vԴ�P�h�{wa}�O��_`� �2�JйR˖e�~g!�$��';�����>c��B6�ǹEi�O��=����C׏L��َ"�X�S@"O�8R"G+
�ܜ��E=���W"O*4�F���:�H�w��2��6�'�!�7kH?4�Zh�#�g��"Q�8��I?9�p����|�3cAݠg����$5�I۟`CקIg�^���DY�^�9�w�'D��竘='q|�BR�����A��'O�=� �����D/'A�l��J��G�H(d"O(Yd䜕
)$���I�M���Q"O��Q7�ɓ_�@pr�H@�#����"O8�I�h�f����@F*M�\K�"Ox�$�"�Р�`�Ev���v�C�O��8Z�"'�0�C%�4���X	�'Q\���N��ځ1�/�<��RN��O>�=�����s��IU,j$��i�����*��I�v3���pE�o*�\�\�B vc���MN���Ĉ"cy��L�}S�����aښ>���9���B���>?��\j�de�X Z8.�Q���On�T��C����@
ƪ8�� N\4%�&��ȓK<�Hå�U.Ț���S*m�X�� A�x�!�<�z��#�Ϥ5�2؅�Kj�0`d�F4V�$\$aS��ȓh�4���%�9i��d`���!D��}�ȓ B��G蟹`�L���!M�`��W��MP5/]*#�IX�Y8vE��y0v�:��-��@�2K� ����L��@�D��"�>,h� E�F��ȓ1�y	p잖:`A X�,���dP=Q`n�o��T��oW3g�f��j�t,�KA�k~���/2Z ńȓExe�Ġ�F{J����)��p��t��m`f�C.4���x��̂@�`�ȓ ;2����}F���dE�wЇȓ;Fl�bW	X$v�Lhx@�1�l��ȓ1�V��D`�;6�З�=W��,�ȓI:xH�,��-��K�
�tՆ�|{�q"3d��Y	Pr�t�A�D�y"+^-Z�x�pG��;G��Q��ya���� �EOܜC�̰k�D7�yBƒ� ��Q�#�17�
=3VFO�y`�'Z@sCT ����D���y�d�	#Y�,Х/ٸf>����5�yr�Ī��1OYZX���'dŜ�y�}����;�$�v���y�`��V:\A��M��.�H� �y"��({���:D�=f�(غ6���y�@B�����,I�
8����)�+�yR�Тd��H�ǜ�mjН�R����yr�	
��A	D���d���2Ŕ��y�J6
����N)Y���"e���y�씇=�9@k^Ll���b� �yR$�"d�l�V �3�<��BC���y2�I�o$����a^>7�2�*���y��Q�_>\Р@� � ���ď)��'���q$N��i���

0��y2e���d�u��D�*���(�yR!�./L���c�f�6)2!��-�y���=i,z�{2��m6lt���ڥ�yB�9h�FE�#!š~����Ȑ�y⋞�A.�Bď�o�p F��0�y�Tg�Ѐ�v�H����v����yrGP;c��ȣW*_��N��C���y��ՠNy�+�
 #*e��"�*�y��L�cfp��Ȕ+�6��A�K��yR�^y�q�K�/~ L�Pe�y�	8"�č��H�w<8g�[�y���5� ,����?�<�;�AQ��y�!B�=ߔT�6*��P�IF����yR��>$t��H(6�*�B5�y£U�+�b��W
/��uj�ğ*�y�i��9�H�-$^�S�bS��y
� �<����=L��mX�d�e rTz�"O`��۔h!0\�ŔQ0�ٓ"Oh�v�9���D�]L���$"O68�S��R�|1�I�!g>F,H�"O�2��Vט}��,��3�"Oб u"�uK�|z�n�]�%"O�D8�n�v��2��� ���2"O U�%.A�\H��HGo��P�
�	T"O��j�#Ҽ2Vv	�T�S?2�\T��"O�����:��m;3���G���s�"O��VFU�>H()���Ƌjq(��"O �paC�@5�$����OD��s"O
]���Q'=jYx��)1)�[�"Oxd��n^'Y���f�#jhka"O�4����hOJ��t%\'�� �"O�Y"BmC#��l���D��&"O8��u��.Yf"5QQk�Nd�xk�"O>,�PŁF���j��\S��
�"O@�Q	��%і�1}��3�"O�y)G�E/5������U;t"Om���m���c�6J� AiA"O�i ������KC�*�.��0�iF\л7�'��`����(#���eN	Z�f<�ד9?`E��6?�0�.6V��Te��H�P
iXB�<�	�0n�J5j��̑��<�Q�NX
!؃�(���ˣ*=|�d�3tm�j���"O�Xg�ӜC�j���O��2�)^v�qO����Y��c��н+� 
 ��1M�Ν��,%D��ӌߑ�!�/,R|� �IE�1��1IA.�O\���oP�)����M�A?U��',�]S��PO~�lʋ>B��# ZD�p���1�y�I."�) �O��m��a�dݵ��'Z:	[W���d�Š\Q��P��Yb`V���J1�y�iʨ�MaUdVy��sQ% ��y� ��;���3�J�E�uIQʚ�y���pHj�ST"�:=Z��/�yb�ǽy����A�3=nͲs�K,�y�_tV�%��@<*��8�*��yB�I�(���jBHտ#�t�e �y�U%�*��5���gž�y��@?S��waDS;b�zD���y���>��|3�GK��|J@Lѯ�y���y򰐊D��a� |j�Q>�y��9:
Tt cO��W؈����#�y�ɍ4tlu[F�ŦK�f�kf�\<�y�_��y��-|dx%�N:�y�m 9A��U#�eu!䥛��y�� �j%XTy2̦d��*�(�yR��X7�t唪X( mB�oϹ�yrK�v�X���.�R��LҖ ��y2ep��ӡC©IC�����U#ڰ<)�c�S���Op��`�_�N�" P�+�ި""O ����A7�%����:mFQ`� [2mš]v܄�Ж>E�4�-^/�=z�J�D��d�4�y�iS5[�Th�խ!w��x�P�^�0]���O
�St`����&>c��{�s��԰s_�J��@�@n)�O$�CboE5!倔�p�ddaD��f���h�!QR@��Ɩ��	���z3��O{"�S���7C�鳰��!��၉��=G�e$�[?�q2��z��ɗ2���j���x�� {ƞ��y��,t=B�כ|��	�)���y��G�B���?R��\Fnt�  U:w�U�(���i��m�'Y�]�O��!���#�I�M�E�'��h��o�:'H2i��I�q�V�qs#R�#���q)@3���!�*T2?.�2���|`�+.G�T7>)ؠ֞?�T���8�)ȶ>�:�����|�o�	Xvh��FִP�	)�o�?K��,e��#|Fraáe������Ԯ3S��)�W��7V�) OJ|��h>� ʨ"�j��:HLcF/�73��s�%3���ڲ�B߀��c���@��@j�٨	>��uHM�BU�wAr��؀cS��R��A�s���h��xC��j���'�Z�W�p�H��O]��A�	z��aU���Hx���l���w�:��Q	A���etdj�
�O(�&n���(D�c\����j�ʬ1�.�0I�5)�`={fa�F�Mg��`Y#��e��pW>�SC���oG����C�u��_�%��0 �K�j$�1B�E�J_���	� "a�� H>m!�9k��l�T�
�ݸ�"�0C�8�)p	 �}�X5� ��j*�4M���铚�Ԏ��$���`Ś�p��		�hO�C��I8ol8qƁ�Xv�R�^9�d�֭@�6%�6�t�R����e�v ��Qf�	F%�Ei�~�*�`$��R&]J�%�3n�s�V]k�k�O�m�D���:��h�(��"��
r�ݗI��=�N�~��(T1��Ȼ�Wg���4cG�e?ֹ��L=~z�	I1r�H��'q�Ա��L�h���aO
:]%c��Ϝ9	Ȍ���	����q�Ѱ�ug'�6���b��-��i��q��$	�\$@A�ŋ���3�G(�O���SĎ;��I��l��`T�q&��h�ܹ0���M�X�31FT3l2���n�J~"�L*a7�L�5����d͘8H�s�m�l. �RG��#UQ������@֒}`�&B�)qr��O;��ƃ�s�$,�b Jî��ZV�	".���v̉-��g�{Ra����E� 4�.�P����t8.B�!H�s�,�����⤹G�$y#�0 ҂��,���P��(/������ʂ /a"�el^�At�!1��P�A�cQ&IQ�6O� B���(���diP�y"ȡ;�'��hb�ʑ<D\���·s������'���BI,};�bpJ
�h[*��Z�R����烊 ��Й�%	+�=�<E�t�Mpa��!Y�Z(ܜ��X��On`�Ы˟���JI~�c�C�KN�M{�iX�8�ԍ�N�L�<�잶��
�I��2����cy2h',��&�,��'�1��� 'R<��,BA�3���`Q"Oڜ��	�l�u�JйY�V	1b��(�$��!q���&�"|�B#Ws&���o�d�T�*1��S�<�G�>}�B2e�هe�!BFky���2�{�lV���gܓF	P,2�aW�#���2w�5�����	�D@��/߃VEABC��.�N�q���%Hu�'�>PY�_	�̂1gX�%��Q{��$ݲ}/xؓ놝`O�`rg�a>E�'I�&��iV/P�f�D�A�*P{� �qr�)�O��)SEJ	޶��E(��V�2ygY�p��"GN����ܤp�\��'-�v"t ,��ɞ
D �m�邬��� 1���!��*��)�Cʫj؁�䝓d	Ҹ���^#m>����f�(/J�)���j�	M�SX��2�aލrda��<����Q��4M?�O�B�!HQ́��
Z	G>��R�E�.��	Q�^��:E*:lY�n*�H�D{�&Y�xN�P#bN�(4 u�Oo�'��-a3mH8JͨP����;�B�Ivh�6�R��|�U�~�("��A7�J�{BNWX�q�n@.b�Xr.T�3�!
b�#?d)~b
�kd���$���e�CEڵ��fA�FC��AVb�p��ԷDOJS�[%<f,B�	�*���&��5�h)�FB�C�6�����Ff(�[S ϗae8�H��C��
�f�4�h!�B�2��*� �s@@�Zn2d�@	�8���!9 @�X�!�O��Jtg���dsS�*5!2Ō�@s�, 0�4&�1�/�&Y�T�OB�'�B�0r� ���)J1n�(�ҍQ`[v�H1�VA?��ʰm�& ��ċ#��#`�[}ŉ�2bn��pb����ɘ��0O��!�i����R�1N�
#�-ט5�VC �<-Ic!D�����-e�e	�H���Lքi��ʼ;�A�$&lb\�� /N߄�jaH�F�' > �P�S�O @����W��]з���R�2��( (�����3��=�*�C(e�&�|5��'���O�h �����m�bɓ9��������M� �>�iݹӐ<\(m
��Խ:W����4.h>xT
�Y��C�^���E�ȓ{D|k�"��{�x��ѥ��>)��^�؂�Ȕ��!�Q�B���K��,����^�d�7 ϕ^6ep�g�5swa}��On����I�U�­�G)��']|4� .�)1�8�k�j]���Xj҅G��ְB�N3����-4��!{���<$͘C�Ԇs<����!,�Hޱ�| �%&S/(�Υ�e@�)�$*+�����o*o=�4h�����8V�~�<��'O�DP&X����&�"�d#���LSDu�'��dж���WH UrAhF3p�g6Av�p
�j%T'�	�+��~�'�	U<"���'L�t��DǬ����ÇzZ��P���B�y�I����%5(���2��h;�/y'D\b�d�-݋�"O�,�d��xҨ�ك"�v�=��Lb�DE+���N@d��C�7���C�� ~ ��0U �#�xţ��'n��3�8>af	�"B18�(R�N3� ���FW"*!��K"W�@=S J�9=db�Ϙ'&�ѩ&� 3�D��脻G�x`Óh�9W�R?����|s�� DIr4n�k��}{�D�x*j��u�T�D�q���6%|a|�-3ux���f��>)�ŊW�Ԅ���|P��_���S$���a'l�� �"�ӣ	�*�I፟�\JG_�!C�C�	�#��T��,��|:�ٸp���R�H��ʅ?�>,�w#ZȼM�l`��v̧���$"Ө\�����3D���	�������U0B��;Z��+5 �&�iJ��N��'&B�4`K��ϸ'��0��`lu�X�% ��Qy��k�H�1+�	8��t���$��-ް �@ �U@F����c��B*=����	�8#.����#��SFo��@���ړ���,�А!*O-[�Oz�4j#�����'�����-K��p�wJR�h��J�'����T,�fs��yG��hF��@�M=J��`�g�t�Z���ψc\P�DD��J��nN+]��z��I��l��
��=!��@��&��4��h�������G���y�R�&�R� ��b�٣U�ϫ��'���zg�&�h�;sZ,	��	�'m�uQ�I�R.,C�ɷay>dKTF@��B�@Q�1�,\K6�´AmX!,O����Y�� R1O&da�cؾ^�.)��M T��UEϕfJ�8@K��v��ѡM�ZP�@Q�A�� ��ͅ�	�{I�@�uK|�F!�v?��dW(��ˁnG��?Qb�>u��X��g�U7�4�N�{�<��*����y���4}T�!�À�\��DsX���՘ǈ���r���T��L�bF>QQ4|Q�*Ot�J$��:ʅ���>�!�	�'b�U�W�eb�
d�?ftH��'�~�`w�x �t�3�ſ%܁�'��݀��g>�e�NA�vM��'I��!��-i�T�Y��Z�E)\a��'�`��$�U�_�*��`�8r4{�'��i�NC�|�f%H��²6�R)�
�'�Xi��U�_ظMA�)G57ﾥ!�'T^T	�[���f�+&�Hr�'���Q�/��N^
��q�� �H\9�'��P���H�L��Q�aP�yJ�:�'���ȑ*,���'��+ H�2�'��Ղ�@`�I��HG($a�'�d q�@��7K
C7TyB�h�f�<�L�91��2f�	��h� �T�<��k�<jVE��'���	w.T[�<q �z0P��]� `a�W�<A��,8��Y����0�`�X�<Y�]�C���+��j[^��g��~�<��"2"�Rըg	�:rt���l�<QG�;P�M��lB�b�L���fMm�<�����5Cu�c�4����cEB�<9�jQ�69椊��f�D��I~�<I%�%y��́�G�'8,�5��W�<�ҍ����.O�y�z@�5ƙH�<!���R��@���θb�@D�<�����rچX��dZ$A%|���B�<��`��c��,:wN�V[Hk�N�z�<9��;���B�,Nqn�;��x�<AGپw�P@P��^y����K
L�<����_>21�D9�6�
$�L�<�)��w<:1��*E�T9��
o�N�<I�A�8��I�A����W�<1F�����rD�T��]R�.d�<��lS�?�B@P�ۈ^����4Gd�<1�㖊6\ȼSA�C���5K�g�<AOΖ^�$h�]+x⁩�c�<QB
�2w�إ��5|w>y`��Z�<I��Z	aT��$ڏI�,�H�EWV�<�4�D*5S���̧P�� ��V�<�� �R%�x�%�u��0��^�<Ѥ��5τ�`�хb��0���W�<� ��ӭ�N��y��� t��d
4"O �qs�+H5D�cGJ�?qz<Y�"Oju땉�_ל��X2h��1(R"O��B�� �����_�ZW��"O@5*�!}n�[��R���\Y�"O���7��ۊ���ɾO�X
F"O�Ѯ�X��](D�l�1��@�<�@ˍ;~�Hp�Y�{Zx)��F�<�Ղ\�<px�+Ծ��X�S�C{�<��m�T@�KG��2K���bř{�<�&�ٳgO@X9�L*'%�=:&gLs�<�2*	k�0	(���<ܹS�FD�<9#腓?b��q�_|O�-�CA t�<yP�>s�<K��5RIV��\�<�'��+�2�a�qNt���O�R�<� �ߵA�L�b�"R�̒�V�<�FȢE�ȼ�q��0��Y2�i�t�<A�F�)�������VY
�!���Z�<��P=F�Խ����7}��`2��y�<1sf�/&�<ҡ�U	�(�i�u�<y2�R)�N|ӗ'ɵ^����Uq�<��Cާw�0\v-��qZ������V�<y��J�&`�$��e.�,�t�Td�<�c��pk^U��N���X�bI�<Q!�-k��$p����H��q+}�<�7��EP&�w,C�n����WbGA�<y��A/P�հ�g�=(g8����M|�<�E�.w��ш�D�8LV�9���{�<i�MY�J�[�G��l��d���Y�<�2��F>�����(�2�	�'Q�<�Qe�=��e�7�`^�5���FP�<��HD������ D&� aKR�<a�E)���rN<K��`&�[O�<	Dl�(�U���B�"�h�#�s�<��ϛ�O�T@���<y�=�"�s�<a��%F����D	�9��r��m�<!r�O;�L���皰�L�C�#�m�<�ÏD2
��ˁ@�T8R-�M�<��ĞX�0��Q�)J��XȆG�S�<����`�����@�X>���U@�<q��)<���rV��h������~�<1��3"��Ս�Ae��p�m�y�<�$N^77^�yE&r��8�Q��x�<�� ս/��y���ȡJ���9�p�<�׀��
Y�y+ҩ�**l��a��[�<AB��5=��P��n(8�"�~�<����,]�1�ܦmP!�a��{�<���	we�	ು�@�)R�Vw�<�qG�r�(A�e��U��P�QCK�<1�<���d��,�Ar�WA�<A�U�W�Ν1��Jb8:�CB�<q&DA�*��E�!!��]˵FF~�<�r�G,�r��\H��KX\�<��׼"����ꜜ:d��Ye�Q`�<a�E�0�|�cU��8"!��f�<�V�� ����`T>s2��!'cc�<��`ŕ^	LI��o!�`�fn	`�<aC�H�X���t�۽H � 2��t�<��!ЫuL��v�ߝ[��� A�Y_�<Q�F[�`ȷ	�
���8w��Z�<����!72P�Q���$��e�d�UU?��"�<���'��b\��?��G�\ wEn}�-��~�B� �*�On��EBE�WJ�ֈudV(c��y/�����\l�D2d8
�ׂ(��*Z8�eSu'R��e��⟄S3ҐW�|�ۆ��*!���� 4�`��N�]Wlī�h�zڨ�Y�X�Ao�#z�}���'a��(�	ՍLK��#.G�]ub�@T&Ȍ7�D���� :�vp���O���rhM�c*̡QM� ,ʦ�Qga3 H�sa&B\H<aT@��n����ʏw�q�E`��ǻxc��H�@ۆ�T�J$ 	 n���>��O����%� V�ܓ(��q�����X�l�z�銝^���[����r�(��A��ZŰ�{&�P�)נ ?,��L;}r��9����l�%$Mލ���4|b4�?�Vcώ C��?MB����TK�,%���d&�%�14��'t�p�d��8]�ڈ�剉}��P!�/F�%*g�V�H�ЉXPǊ���d!� q�j�D=�S����cq���g��1�G66t�H�C<[��	[��'Ò!8W�G?a��	1������3��g�z������K����<�H�S�G>g��	�}�v>����,#�l�i@`���{"+6�bl�7#σ[��G�[��U9��ҹT�$!�0�ܾg9�LJC:�<�kei�6��[�#�%5�T����O�����B��Xή]ip��K�Kߑ���Y5) -�b�|�3���d��J�IN����1;`��+.��툥�H�z]�es7$ �M����-\Ο0����6vBaz�#�Npy{5��&/6|��@�����[�c 4u�a+F.�0�mZ�MfQCE�%)9n���ueR��dx����:��6JQ��p?AD��O�J<Cf�_n"�H��$�j՚��J�g��7�Ļ�v�pD/X���?� ��ޭ[��ɍXX�EiY/\(�%W���>��EQ�]��])��%�S7^|@�����ZU�uDU:O�h��Oĩ��I(q��%>c��)�JؒO�>���NӬ~A�bϩ�t��	]�q�r��Л>�}����PȮT���66Ȋ�9���~���@$���J�*`��	�`���j��I�I����	=���'�T�y5E�$&|E�ɚ[
� �c���ē4�@\q�ڙp���rT���O/����>�p�:%�rs0dZ��(m��dz��ʿxA@5'c������e��b�"|jր��jN0M�s'Җo':�J��j�'��D[�Ɋ�:�q��4���+y.-3��3�����"O�0���X�h���&�["C�Ҕ�Z������n��'XN���H�',}�����'S���P#Vy<��ȓy��qH��p��#l�e����'"��ja�؅0�ɧ�ʹ������$uA����a�aJ�"OԼ��F	�-皴8	�7a`Y��{���u�Pr\�ϸ'{����!	�.W��y���"��Ya
�'������:��0󓈌 >�l$����� �S�,�O�գ ��t�Mђ�
�(D�D�	�UWƁ3��)�F� �S�|�A샢F}x��2#�`�T��z����a~$Y6O�n�c�8
}�|��@�Z#剣bH<�y2M^� �b� ¬'�
��"���+(��X(�/��}Ɇ�U僴b���"O�@��"JÊ-0�ˇ�@%��*�"'�05�d��rPj��D(���|툴(��W�Z� A�f,r"��!�2�'m��n=����B�r�ڀ�!t*r���0�"Lb�릟�1��C����7�"Y=xE��I�{�'z�Cec�,9���S�"����$��H�V�̢I�V��pB�_�TћS+Q�]#�qqG�Pd7@�[G���*��V
oY���dֆ/u Q�A�Gp�3
��P��I88�&�%Q��eXe�ׅ*r
Y�a�\Bn�ce�G��ѶQz�Ek�Fب}�L䳄�I��y�+��C����V
�wݔ�p$�a�|�[:i� c��	@N.�8�k矈��vJ�0wݖ�`$dC�y���|Zh0�p��3��yDO�0>�`F��p}����7nx��M�!�ʝK@�l58�"C����t@"�]�f`��6���?��p�!���a���p�T��.u\�$#�eN�<E�Q���O\�v�Y�-sV��J�*О���BIY,�`c�t͂bY93"���G����nV���߁yV�UZ���[�v���^�ȣ�L�"Q@����w����������weU��$�{R`Isg@){���	�'�.x�������siK��d��"T�m������n6E���R�B��W�	�!��'���O���.I�
�F�8�;<^����'HD�f�Őq0v��b^�]�`7�@<!,��+5,�,(H! �6�!򤃧z��p��`��`�a�/g��I".5�a�gBAW��e� 韹2�>�ҕ+۳�Z���TSp\h�V�>D���mF��%��ES����Jب+�t�����Y2<�a���x����qO�܂❼y�����F.q��%�'�����b��X<� xĮIl�b���a���)۵#H�D���jj؞�iC�
FN$-�@ϕ�~��1V�"���e��'����/޽5â\��'j�	>�O2�(�N�F!�DO�����Rz� a���
�	�v\١'BE�0 ��F�k�O�x�s�B�W�^����,���� �!���'��L�u�$k(d]PEG�Z���J�D�� J.��$�D�"�K��8zL��aAC�"dV�G�f��DE��v�-���Y�,���*KQM��I
��L�F i��y�`G\�{U���D.5\��;�DT*zd�	��}� � �mАX��$m͊E!�ߢh*��&��I�D�2\�E���ڔ&1V��s�l�X�mĈ'y!���
M	����
�&��"%ދ2�b�P�a�nA���'�8,ڃ%͂S�y3�B8 ��Ţۓo$
E W�T�Z�R�䆞p��<y爞���TN ��!�$�4-Ԍ�6"�,�U.ٞ�qOp����X��q�F�?�'R.`��B
4M5 &nB�eT��ȓp����T��#!t|�+� A�w�RYK�܎J�$2bW��k�<Ѳ�R� ������.-�ؠ��p�<�FG�*e�h���E�$+>��(f�1ivδf�oR�T���'ed�2fO/#�^�sԨ�,�X�B	ד���K�%�^���4YEd(3s��8g�,���J��܆�!Y5�"�J-��zc��=A>��=!�"\9�H�H� @���U�/m� ���C�;���F"O�y�2j˽J���"�"�"a�K.�����!zy�-�m���-d,I�w*3y�4�a��f�!�W_}�T�&k�xS�<F�	�t�x���G�$n��L�gE�S؞��^	J_,�y&F� y
0��D=lO�@1�����[��=A2f��f�0�r��>ax��ȓ;�Tu��O�0�x��K�R]�?YV	ԪJu����	�}Y��*��T�E��Pӣ�#&*!�_:>��;���x4Q�ݫ~!򄅿4��哵bӮ����EƱW�!�D���D�t���|Hy���*�!�RTx<i�(��U���tƔ/(�!�DM�^lN��G	J��8�'�+U�!�"9���ӏP/i �+煔27(!��T�1����
E��ع��>6e!��Y��(	�&�8�,��"#�%U!�dI(��+��ߝ	��e{�`��V�!�ĳ`8�X�	Lf�hiI����]�!��|k@X�c��*�v�2�-�!�d�<iѴ(#e柝t�BQ�'N�1�!�$��[�IVn܊�x�Η�3h!��-,td��"�۶��TAWlD7M!�$U1t`f�hĭB�O��\��M%:!�D��t�^�[��B�*# h��;>�!�Ą�W�0=�ҬŽ=�Ȑ�G�C�!򤗉c�p����{�*��Ug�&,!���$$Y�do�9e�(��b��7�!�D_�+$L Z�cO&�B����[�!��� �a7��n�aP�p�"O��QC�4t�$
Ů��
`ʷ"O���Q%Me��5FޭP5~�f"O�L32�]<0�ʕ3���/L&e��"O`���b\�R� �r�n�/	3�D"On!���RW��-��q�:��"OJ�yF�F�g�\��2�Y��P`""OT4R��˔b6�6Bƚc��m�""O(`bD�aA�d��N4^�����"O���cՒIZA�P�J���˰�(x��۬<?J	pd�7{�'>�A(r����B�Ic�u����C���*7��a�T>����ێM3���N�(>�,Dx����;�I3z��D�2���heb�1d@�wk.(H�OfD�gKXn~�哢P�^�17A߼eD�QtO�G��7Ͷ��SFaD�����#u�@ם�47�M��D�T����J�p�$L��O.)�)�'�l#���&[7��S��E]��p���ܲ��'?%>O�y:~q���80��r㏏+���Wg�I�W���>��`�*:B[�/��W ���9�MQe��ܱ`�Oa�� D��Iˁ%T`�@T���-k��i�qO�)�S�O���c��aq *Z���3];�c���h�t��g}����"�UK'N0���dh���֮N�bP�{���8<�|ٻ�b�L�8�Q�&D����=;*4�Ɍ{��i��־=z0�	�&�\0(��o���p͛#��I Y��=�)��c�	F��0�(�LԂ5�Y��b	FxJ|�1C��ۧj�D��I �R≪�#<�~�"J��{ L� 	1��c��s}AJ��O�>�qNH�DZ�:�,|�>�g�e���&�i��D���~��D�?��#�G�Kff�ʧ���S��{2b��>c�	�m����D�p>u�*T�Ist���&qb%�<i4푑�@0�ԩ�|��0E\a�%��*�z���S�w=��I�YS������
}1�S�O�\J���DQ��{d�m���� d)rM��L�%~B��S>[ZH�0��$}Z8(V�dSZH� ���}[��C�A�a�t���(E�Ջ%,�	/���O�P��BD}?q���?y���O���?1��LU�mLB́�߁p�L�7-\�o�V�m(9���3 �C	�����(`��fɛ]��)['�D�v���	�K�n�go��a&(��剛J<��t�%q���To�<e��B�I1X������ºT�h���^H	�B䉸>����3+-$�Z�&0Y^lC�	(CBi�#�6[u���fÚ�#�VC�	�S��B
^�����l��?�B�ɦe��YC�kB�t%�q�4EM+��C䉸e��*��ån�R܁``�=iZB��iG
�ѣ�	�ts���y4�C�I.a�QH1�4%
l��#�t�B�I�'|����m�)ږ��Q��C�I
G�`�'�ne	�+ǱK�pC�QH4��� �2%J3M�dPC�I�Vg�`����\�Pq#��)��B䉖>�z0@���
VO�}S@bܱG�2C䉅3�����,��-�����6	6B�	*�f�2ff�N1��(��.�B�I_��ƊD��)�� �B�I���� 3c٦eE�p��EQ�8B��)W]����EB�!����g͑*-2B�	�$S(�����x�x��N��C䉼(�ԀB�I�FV�kW
$5 C�	1=�u+�M_�D�K��Ƹx�B�+>�J���dا��J"�Ǹ&�B��$,�z [(�k��]09P\�XA*D����xG�2��
?�����'D��B�oޠb!�1�/mL��G"D�� 6"�&�H���*նq�&�jR� D�"��ڲgiZp���bm��9�$1D��钇
|�.�JPA�~���cE1D�H7�Vtv��-�"E5� �M0D��z�K":6$�V�_�7���ZD�+D����-ƫ,�>p�n��4�P��=D��$ŉh�f���,Vt��@0��=D�tK��R�M���`�El̔i3�:D�TID�T-r�)ꤤ�rhY��6D���5A[!���q��T�~�P��4D��.��,z\u��4\�ؑ��1D��*����m��V4�A�.D������7td�ن�/�,�A.D��H��Q�k�2��s�@�yiB���?D������&6�t���\��Π8S%1D�\:4��<A��%�P�}d�p(a	.D��B��r����Ę<N��9s�?D��@���>jԌ�#	L�y�9�:D����,t�x4��U��	=D��BW�A�2�r0p��K
vh����8D��kfa}�pۗ��%��ĉ'7D�� � ؑ��L�d��7!J+L7�}C"O6�J����|m�Q�ߊa�`�hT"O*�����=b��2N���B"O`��Q�L=A�X!�L��*t�]��'�A
���n�V9�ek>.�ą�
�'ܮ���/��h.>-�� ��]��'���J��I�*��e�	�.�`%(��-5 �^
Ha���C2QvEB�'h��U?$���`%n@�Y�D��
�'�h�2�P6zt����&�J	6M�
�'�LL��E/��-X�C�P�8��'��{��P�|z4X83gH��p}��'���{pm�5*x�j�`I�X�����'@���6��;uae�HHN��ȉ�'���1�ёx����=B����'��W�o}l�T+��.��!	�'V�lڤ1s��@�
�>�,Da�'H����	ãY��*Aʎ�p���'8�� �Β"`6�Ґ.̑��a�'�p�ш.���Æ�״4��'P�A��V�V@�D��"}����'P�w�^'F�.�!���Y����'�}cEjϦ6k�qI k��L����'��A0s��,ڼ��dB�znR�Z�'��󕈏C;ba���Ĥ\�m

�'�p;v2�Έ�"��<�i
�'Y,�CҬUdV�`�ݭM����	�'�tX��.��y�@�"Y�V4����'�j,�&�B?6���'OK�����'���s� +0舡0nH�H�:�'I�hj'��S������>�(�!�'��X"�
�X���� M�ę�'r��0h�+�I�E�""8���'Oй����4}5�p�i�������'���;Ҭ�9K�J�n����	�'H�]H7�R�8���Qd��u���'d�(��Հ;D�eX�a^�b�:0��'��8�`GM=j\�	×�Py2��	�'PЁڳ/.	���C�C�>�p�'�Ԍ���
HUu��?�0���'���wo�1^�8��
"4�:%1�'C6Y)A% �(�i(���1k<0Y�'}�,�0g��IY
�"4`N�Q%x��'���HD)Ȓ��SE�N���
�'l~q�p�R�<L��f�@�@	�'-|D)�M�L+@9�28kV���'�� y�c
��b�Qa_�X��9(�'�J�٠BIh=쀘��Fh>Z�x�'�*\y�+M%����N�_�D� �'P��������IX�X��$��'}8��tO�9?܎�xF_��\�c�'�}�Q�Q+��8V
��kQ�'ܦـ�P�wX$�P�����p�'���!�H?E��y���H�w��
�'�XY[���*d��9��/jZB	�'��m3�֏W6�D�f�ya�	�
�'�eX��1��ɉ�j �Gg��'�,(��1\�
Q�ȧ@�n��'��K�%Q5��бg��?�Y�'	�և; 3Ј!��ƀ=�)�'����Ç��!��LP�l�^�:�'؆�ےEB�{V���a��d���
�'@@�!�ધjH�(�^���'�V �����'�bm��P*	������ ���Ǝ�0����<���"Oԙat��B�,�:�� 1h��e"O���M��%��t���)�}Ӷ"O���r�[
�<s5d�6z	B�c"O�<á���)P <��E��Z�i�"O�Vc�AE�|�U�G�`hj�"OV���ʎYHib`DU�t�N=�"O  �SO[������ �-y��|(�"O��0���;�m�``�x�~%��"O�$P���GF���ϖ6<@�\��"O�<���sevA�����
��I��y2o��GYF��Ċ��Bq���y�e[=�fِ*�-\�ڨ���ֺ�yrn�Yݾ����@3f�A�,�y⋃�T,%����@D�����	��y�J��@ȸ4�AHȂD���÷b�/�y҇%"���s�E M�l�5F�y����PY6����?CD�5���3�y��Ľ\2<���� "5���;E����y2k��WsD�#��ͣ0i�	Ѕ�8�y��).~���h�	}�\$����y�f�*�j�	W��q���!�ԟ�y�I�[�ZhH��p������Q�y����=�Bd�	o�p�#�ǎ�yBϒMK�򍛸1�8ۢ����y�.V9��ū����rƚ�yRE� :w��j
2m�h�c[��ybA�9Y�n�x߸ޝ��N�-�y� _@�	S�,H�Q�����=�yҊ�g:R� ��8Ek�Uj��y�Ͱ){�p5O't1ƭ�s���y�.��g� �P��1�h��$�y2�#H�V�Ȥ���T���#�y��I5��q��ĄH��]��y�OG�O@���o�w�A���yr
��I?��Ċ�vP�؁��%�y��B�E�����q�Na�q.׳�y`�$&��r`��:�:0��D̊�yr%��;�TP��ӗI ١Q�ނ�y2��	 $| ��%�?&p�!A�O��y�cO�[?`8���T�*SK��y"l�*�|A(�"Y�x�l�P�$��y҆mINd�S��>x)"S!��yr.��Ɓ2bn�)iM>M@�oſ�y�Ȋ�5���1Nѫ6ƪ������y�^L)�%�@�X��R�H�+�y����/4��p�X�M����dj��yBA��� l>	�y�e����y�ƙO3�x��l��1吅3U�<�ym�r����wA�%���ԭ�0�y�AP�2��6!�($��������yr$�F�T2���%��a`���y�̉�J�D;_e�9�	�`�B�	�hN�&M\<O�����H�aC�Ʉ%���u�SRy�yIqgH�(�B�!eBLA�ϊ�fVmc(�"]�\B䉷R��q�������,�*z"B�I�@�6��'�I2���<V"B�I(S=�h�vH�>_��RVaҽ��C䉤q�l8eO|����2L�?��C�	$*��@�ŊWL��k��$�C�ɖHi���5M�/�ހ@E���@�vC�Ȳ��2D�	�͸�˲=-C�	*�&1gi�,�<QA��
�ܡ�� ��� �+2r��XG�NO�̙��"O�t�O�%����ǖ#@�j�#'"OziPf#ȗKp��e&��^�\��0"O�b���#w�>ݸ外!B�L�s"O����\�k �z��/�$��"O���%�xp|���/ۜ4iޕ	�"O��A�ӎK"d��%؛Z�`q6"OVH`%�d��Pcd��xX6H9A"O�YĄ� ���
BOd�e"O�IPdn���@�B��q5�Y�"O��J�/�u�(p���Av �"O8`�w���Zf��(^�%N�a"O��#�Ntk�\q���/�4�c"O��z�JG�k�H��$�\k��h�%"O�����t����dM�2���%"O4�@#�Ȭ-�j��aڿ�,e�F"OZ�c��I;2ɪm鳀-	k�TaU"O�U�����	i�b�OU0hK��"O�U:�/�]��1�lV�%g�-H�"O���R���xg�����Ģ�.�C@"O$|��(C�XqP�=��4�"O�T    �