MPQ    x    h�  h                                                                                 �gI=��	�#�V�)Qv�@>A?<#�Q��� oс֬9�`��v\h�2�`aՀX�G��u�г�,�6k�M3ɗɥ���
�m����A�bꆜ�S�$M�z�k�ws����s0�z������a��@Yޠ�{ch�N�}�
!X�9	e�ɱ*��D�q���+A#����oǸ�c[E���y�:̿�vp��%Fs3C��+{���ݺ;+���g��^V[�B9Fy1�_�Sn	�& @��Ag�EXɯ�~g;�yIbi2ܒ�TX��G=���$��)��q(N��-�G�_��S��a�����?<�3��X�	��+�nc��G��j\f���?�~?�0�!7����0v��B�} .s��G����4�&���͍(�!��+�|�d}���2񜮱I������%� �/��,)���E����_�w�@��ˌz��$G���U�г�X;ho,R�¡�������S��~Y+��eE'�x�t%W��D����J�MO�۾������j�X2�(|b7լ;� ����p�d����c�fϦP'-���7GS����M��3%��uԡ��f�X@b=.�#P��wL��k��aə%L�}*���%���B�q�������V�匐<�2w��T��k���%}���z�r��)�xl[]U�{�:����9��(�1�$+���V��q�i����P^��6^I���犪���U��ڲ���qOj��S̗Ut����j�J�����E�5=\S}�f��Ct�iv ����W"k�WRIg�&A��@cW��6+@��h�!T��qiwN%�Y�z%�ީh��WX�\��v~-8����b�"�ʸ^I�-u�+h�Oc��;Z��v�P�BC2`}!�=�O;�!��]x�:{�ǃǗ`�AO�1�|L�I!�@�m�/N*?���o��>����k6w�$�[V�;`{�!���< p��*g��1��r��%���n�y�h��COVoW�'� 	�P���vnBx4L��ef^C�ׄ��˓�$F��-"�$�L�U�t��Ku2	6�h8̄�hJ�-�|х���俧�7h�xzў��ǁ�GVft�Ê;���&t�w���s�Qu�='ˢ���6W�k��V��H?��,1�XV��PMK5�`��\E��˷ϳ�Jr��D�Òi\�Ҥ�RBb��S��]ɻץNo���LY�ȟI0�_���x���/Ct���s����m<;�cN��yt�%l�H8إ34����Iu�A�y�����n�*���Y�{)�k�⯏�q�?�$چ�Z@Y�uTf����e��F�|�Z�}�:�ET��cv^n��t��6���{�ѥY��QQ[s` ?FV5�<�1�s�ς�����?il����k x%g�w�ř�=w"a��2ɷn��t�;���s]v������g��䁿�S��s1�tt)�g=K�d$ɹ���	'2��"�_{�A���԰�P�A?��?�z*�s�9����
n��FLٌ���*8K��w������*^�P�+/XT	�	i��#Ng���YӲU�5��O����7}������H(�|���uce��vk0�����P}���1���#aL�?���+�'ۄ�H�8ٛ}t���}����չ�dnW������"�o�h�C �S���MT^�ł��g�~��)Z��}�����'���b�]�l-p{�l��ۚ"���!��+��[�����|b�M�B�/.��瘛�o��\Ps�x^��Z6=%M�m���]?$o���\�"}C_Z�L�/ӄ�h5�2�H��D�~�\}6��ԏ�ÿī�c�~��w:8cli��m�!��&��Ĩ4@���c5џ����M�u�����j�Y���U��Vs���"�O2o� [^H�LK�&�i��aacMԃ���V�_��v�A�\8߳�͗�R�y!Y�8���Vp�w�V��Mֱ��Y��B�=~�_�-�XK���tN咹����B�Ҳ�c��A���9��[,[�.���� 3�=|���o��{Q�cl�7��`Q��OD�z�g�W%��� t*�VA��3>|#-��[v~�����Z����`9;҃J��$�9�3����m�b����YiLG0�)�_�?gL8Tr�'��Å�%��5/ş���� R.5�ݒޔ��\�3,G@�l�¨�����G��*����r�#��޲ܻ�+�.�ed�g��<j�
h�ՔO�g_iV��]�
��q��wfrR��u��%������l�>m�܎�z�?|��&띚������22��D$�ȵ�r��\�Q��?����--��Llgt��q$�u�"5�����O%�O��ާRT�j�ëUi���jEfOBXEaT�
�Ïs��!����,��'����JՃ�yE9�����f��i�7D�'��;g��3�4�X�'��zX�l����e�y���$�}����I0��W,�H���FyVR�q��ӓ�{�f�0"�HQA�-��g�Gє�����m���Fׇi%��3~�]U�}���R��ix0=b�$[C@�S({��Yf�jDǸs���Q�uI��@k�a�>:�����V)E�ǃZ���a�D���޴p��G_�(�t��5�S�בu�*�0:fVjw�I3�&k1Y��+o��)�r�SK�T�)ؒ�!�GC��/p\ҏ$QȊ�
~mW�W9(e��&H��7}÷���9��p�+n�x>Kf��y8�Q��C����Eθ�l����#�aE%B{�i�c�S�Λ����d��w��l/m&:͟��V�� H"�m��k�W�e�/{�HR��w���ڮ}b����Q��1|��w��y`�Y��M���,��o���iHO0E��D�y��|�$+��ۆ�UGEg�����l_Fh���y(�L�.��n�~�f��YUE�he�Ad/ w��.@�ֶϩQ� �@��A2mZ��
��XC'�8�X�u�.àT�1��ՒK�V���l��p_37=���)�Y��uYZ��!Q4����-�Y�@9��<~Fw�E�;�r�Q��;��v�S_2��@a�&C�u�1�ڔ����M,Fbި(Ρ����0�]m�'Q<��b�"��n��M	��k̽����L��`7I�<g�>�3a��9YYb�{>Y�N��L
���9lW�$�Ώd��q�n��M7��%o��͡a�E����B�%:���v��"%��]CΠ{���U���X��3�y[x
�9]1i8SI��&[m���;�@�ׯ�sYg�H�I}����X�0�GxV�ѤNy�Q�qO�N�`����:�S"ܲ�&���^Ě�(3�5-��]	�K+\a%�ȕ��rp郻c���d?�$:!Rb��}��0Q�>��}����۪�h��b�T&�B��H���;�+@���h�ؑn�	�7�����w#��>��6&�����_a[�2!q�.���a����E�U$���S0�o��A�\�S��­����Jf;�e�Sx���t���U����`�Ȕ�ۙٗ��hjo�a�#�70�������^�du)��>{.����-�ʥ��FG���^�N������Y�ۓ�6=�d�P�L�绯���@̑�P����B�dB�h�q��#|Ǎ�:� ;<����Fx��'fN˴}����rh5k���]���{u�0�ɮ{�3k(䳦$�St���q��i0����^����&�I�X���G͐��!$�i}�L�!��>��P�Uo���qJz�v���G5�� SX羋,��X �w���;k{�I�@�Ap�c2�+6f3u�I�!O5P�̊�w	>,Y�-�$�h�y�W��ŵ�<-3))�R��"�n�^5d!��2+CcM��ųk0��ԫpgC�:!/�w;u�rTʢ��������O�Ǣ1�mu��5�@z�/�I��H&��H��r����6���Ey6�+;��ڝ���7���Jojga���9���t�|��m���>��o�R�'��	��ll��ɮe��ҿ��e��+4�ʰ��2��02��?uͻ��c> ��-�����Ѡ=��_K�c�W��zl���RG�VZ�~���JtN_��4@ߌ�+=�S0��%uW?���x��c����Rس3Sl�N1M�(�`�NG\�D(�r��e�[����me7��R���N�p�:�`�8�5�L�r��z�J�����؍�,/�(�K-�����m�=@�>��ô@%�8�m�4WK0���2K�y'ě��n˞w*V�bY���Ɩ��Jɓ�Z��$�r/�5������[��e~-�JZ��r�Ux�EϋzcQ�U�"5F�/��4,ک{�%�Y��Q��s;�F��E���1~g<��S�<��i�k�[��x���g�;P�4a�=r�G�s��2�2Jnڰ���b;lGs�Ee�`���b9Q�܈oS@�E1� �)w_K��_���_2I	"�T��o_6P�A���+ceP��?�l��n���
)��Fg;0���<K����Y��j���+��	�Vn��s#)g^�4U ����+#k78)�����p(�'x"#bu�20�q�p�i&������F��l#�]܅ڼ�a�������O���݆��7��A"��{OWR��B��=�J���} q�0�W�5M�l~�}d�g�̺�5����~����}��)��]#�Kpv��laEK�U�����A��_��6 ���Ub*2�=��/�3S�S��Ɋt�\�q�S�Ǖ~�%��I����?��NJ�=�s}��ϛ'KNӿ	R5t�H�DHdk�����d�>S̫�f�~�H�:ӈ�i�(��ǿm*���#4��u�>�!��SC��z7u�1aj�~���y�U��sjlի]S��j� V��7�T��
�i��a��4�d�FV�����A͖d������y<�7�E��1�w)���~3MѶ��<B:ܪ~���-Vc�K�y��
��-�����a�-��c�ЦA��
9�C�[`�.�i��<�>����]�!o���Q�`��}�`,W�OE��r%��[&���7V\u.�)�#�[����'�U#��,��;��o�|�6p�3�"G�� ����|	鏴�G��J)����8/#�'ݑ5�yq�0�ڟ
h��Er�.!ޚ����b��3gl��i��q�3��oϕ��h����@e����|�ƿ�`�hg�
%��e��v:1�B�9]<���l��w�����ڀ�X��u����%��m�܉�uu�|BG��X8�����*7�,���0r��>�L�?zM �fVD���Hl�7�L�%װ��5e���qXO�S�q̿��}���>��0�����E��X�TY�u�J��<�v�u腻⢼�!&Jp/�y@&��7ϰ0e���DL��g���&���5��A�'G-ez�߶���e]���X.���3�I&0���,xL�Dմyq)�qE�8����fGD�"Q�mQ<�_��<X�h�*sۘ��@��uE���}]P�r��IR��V��%#=��l[f�������a����sF96Q��I�k�l�>uc�9׺)@����Z�\�a�Ǟ�Y�Lp���_*T�$`5������*o��fq�e�13���kl�dͳ.y�t����KPvp)��!��`C[����%�*|�L
�e�8W�E�9C�ȗ��H�O�7�U!�X��ǯ�j$)͆>f�W��J/,U�CRT'�T�����Ѵ�#b$�@\/��=U>�v��v �#w&�_d�w���/(t��F��J� #��N��m�*S�{�򇲴���S�c��Ō�x�f@��}�K����E�C���{��ٔ���"��()��.WĂ$`F�{m�O��n�3��RB|�a�e����)FE����q_�%����g�2�,Ci�YT�59�U�Ah`�7d��ӝ3��R��
��t�|�Z-�%����'*����IJ�Ti��аLʿ���c	��k��7�(Ǌ�D��t��u�������3�!-ga�@4�V<٠ ����V	܁̍���v�^62>\�a��	��1ѷ��1�$�,��=���?� �˥�m����b`�e���M��k�#��9�(���0��&LañZY�C�{j�N0�O
W�=9�����2���q�wS!z��^�}o��<��E{�5睼k:BY�v���%<B�CZ5{G:��.h��C���[3� 98��1��S$�&����w0�;H��6�Tg��.I��܈�PX��ZG�����0�����n�,M.N����׶�S]?Ƶ���߷�����3u�e�8�	���+7tW����r�~������?K8a!m����0,F�y�}6O����^��0��R�&��f���"�פ+{�W��tĠ�(�dN!�#0�9G����R7l�y*Ȓќ���?=_��n�Յ�I?��p1�����F�)U�s��NEo⚚� ��,&���Cˢ2L��e{�"xϸKt�������Ƨ�C�-�t�f���j
�I��c7��c�,�.k�d����;F���-P6ѥ�Y2G	E����i�I�k�m�uĬ�ά=d��P�G�LZe�j�[� �s�y��1&�}n�BKa�qz��b��H�é	�<x5���L����.|}�e<8�Br#�p���~]K�;{P�8���U>(�U�$�45����q��ei��W�Ҙ�^���`�I�{��@�1�e���&�ѐ'���y݉�4Uj �n�GJ5����53b�S3TG�B4l�Mhl �z��o��k6�I���A��c��6�FA��=a!Jn�'�w�v�Y��e�h�<�W�ܢ�2"�-.��ϭ�"O2^P��#��+�vc���N��O��T,C�ݛ!J>�3a;P3�?���=�p���g���O��X1��?j�@U��/Ĉύ�LJ�BΧ�M�p�6�������;�W�A�2jI���m"Q�� A񂚟����rt�����9Oo�P'`}�	��� ���)�e�����C �Қ1�������,=�uh�	�^d�L�{ѻ�u���l��}���D
z�I��CnGg��9��3�ut�D������W!=]�յ���W��E����~.�"�ֳ�2뉟�M�<�`��/\��!�-<��$H�:��H��H�Rx?��I7��R���PW5LOJ��U�U�ժ�&����//�̠�u���8um2`�����%�8�8�U�4�2᣿��Muy�xQ��8�nW*�Z�Y����!�j�'��u��$+��� �����ey��`�\ZH�̖px]EJ��c,$��]����}qB�{Y�rY"pOQ�ws<�F��'r�1y{��8�����?i�A���~�x�|4g	 ����V=m�j��y<2���n�q�j��;G�cs�4��z��]�t�7rS���1���)���K�#��u��s 	��W+_���AיԦ�|P��?/r띰c�i3��ELJ
��hF��{��v�j�pKQ�ɭ4�~�� 2�Zm+���	��;
��#�;�op��������_~ �7�i�T&�~��(q�x]I|u� ��l�������=�����^^��#׎j�u6��͔ݑ~W�5��Lzّ@����?�M��$��|�lW�����\�Xn�^ L�~�==M��n�xf|gKႺ�����-��	����R�d��]��pq�l�������q�!2��"h�3mAb�6f�8/������ɥN�\F,�.�w���W%�lޝ�V�?��*�	XZ�X|�}9�ü��|�5��H���D�Q��Ҏ���#������:~!�`:n�pi��o#��(N���)46�6����=��+�u��"qV�j{-;� �U�	}sE姫���h�5 Q\��	��D�iǃ�aYV�?ͅV~d�A����i��J��yW�.%ʈ�wd��ՌpIM�۱�gB�+~�͘-э�K���>����R��̴�q�cn��A��9��[�`.*F�׏��9����otc�Q�},�->�`'�O�����e%��ZǶk(w�
Vw}_)54#�D[��1�|�Pt�̇!0;H[�o����3�H)c'�
�w%M��{G��%))�Z�5��8
�w'~[���T�+�,�e.B� ].<��݈�n�=4�3�l��uh��2L����*����h�@���(�1�a	a�[>ggn���)�۔E���}�~]�S��g(�w��ʒ�	㨵�L�Ӡ�}`�jm�<�p��|�������*d>�(CE��Sg�>�&r2���Gv?���!���/-l]��'������5 ����O��,������`풫Ez�%@�E��X�T��
�J�W��������\LJ�y;eD�K�k���D}�1�B�Z�a4�1l(��Kp'�v�z�S7���e��~�'�� ]%�z0�X�,ӑO���&y� �q��)����f��?"��+Q7��ﺵ.���?�,J���Иe�ڇ���iM�]KT$�p�(Rx�����=XO�[��4������\����s�Q���I���k[��>��N��$);���9{�<-a�jN����p�i_e����5�ˇ�G��**~-f�f��@F3|�k�q��NR�����(jFK��)e�!x` C6����
�Gl�����Wy�9^���EH�&�7����JZ�&7�$�>���o}6׏C�ť�����Ӵ_�E#�[���_�8���#?٪�F��Z'�wO�4/���\�L� ��$���mDe��vg���ڥL�~���e��{v:}����-6����6_8ٯ���O���W�i@���p�v��O�k�UB��8�|�W��@mF�&�E����껲_�䃲o���^~��7/�4؟�p8�UI��h[D�d���XX����GJ��>@��&Z� ���B�'�A����V�d�T�&�Ћ&Y�� c��L�f�7�w��AƏ�@uO�6��:��n�~-��@/�|<4
���2�q��G����"�v�a2��a�Ҭ�+�зP&�!�b,<���c��z���f�m�i��R�b���� �M�=hk����t3i�M	����a��YOE\{��^Nk
�r�9�ّ���V�ڹiq���C�9��o0m�׾�Ev�����:�ըv���%���C5�[{��݋�:���j��s�[���9S�1_��S�>�&�'��E{6�ȯ��pglN�I��"��PX��`G�&_�P��
��A��jN����vP^�
�S��-�\�_���,�P��30g���	wl2+���>��;�l�y��P�?l!���s�[0$����}����c.��t���&O�>:b�-3+�=Ӎ5���ί����zm	�T���,-kִ�U�l3�ũ�_����~�d�͌� XzaS����UZu��Iz*o=o���_6�G}��/�}�]ܥOe�xʸTt6���ˤ&��鄹�\�O#f�2��j��}�7��W�Q���I�ydk������W�V-�x�����Gd�����ք��Ƶ�PO��	�<=��HPΨ1L��]�%���v�}���v�zgІ�_�B�y�qu���YK���6��<��[�w�ϧ5 ���{}�\,��1r�X:�ɗ|]ƙ�{+~�?�{��h(�\$<6֓��q�Li&?���x^F�g/�XI�U������+`��n��b����$�gUeX���>J�2Ն�r5�?�S���}\6��{ ����~.k�`�I�*�Af�8c���6�ya�؇!E�g����w�"Y(k��٘h��W	���'-){`���"
�^k���P+�bc�h���,%�	ӟ�aW�CcL�!e�T�j;+l�z�(��l?���q��OI��1-��ĺ�j@0��/��Ս~��\�O���+�86�C�d��;Z-��GR�-Op� Xq�`��(7���VvР�菢9��4��oh��'�	:�=�b����9��We7���ȕ�����UW�-e&�����1dg�$u�7�Y������^6��֭A�U±�ȸc��گz�W���T�Gg����ݳ�NH�t[��}�����=�ē���FW�����p晹���� ��T���KMpQ`�|T\V1���d&���|���L�#�]��j�R�.�D��n}n�քx�k�L�A1�0�P�mI�� ��lR/T����#���m��N�����*|{%=�d8�]�4:��z�ށh�8y���uenA/�*�:Yؔ��|ێ�������$���|�&���et:��4�ZՊ����EŲTc�t���E�e�}��ʠ{-�Y={Q�<s�y�F��M1t��ϓI����5i�7j�Q8�x�eDgD$��jX=h���)X{2Mf�nS��;"&PsD�Ֆq��X���{�S���1y�)��Kdb`շAڕ�o	�O��_�_��qA�P!�!x Py�&?j�ߝK0\d����(
�(F�_o�\@E��K����(\��K��a�v+`y8	�P���5#��h���V�&D#���pٵ7���/���Z(L����
u4.��gN��)���72V%�<%��ox�#������Yɔ8��MD��W�R��a?�Έ4����c�w	�W���g�sAل�x� '���ͤM%��s��g�B�Z�����t� â����Y�]Y9�plm�l>���	����)��$���c`�n�Ab`[v�3�&/?����#��H3\�iq�	ŕ�o3%�*����?5�ْą��sa�}����Z{�5!5�¼H� *D�^e��G����H�4ڟ��~\e�:	4�i���~(���S�z?4�����s�Q�����u�� ̹�j6�!� �XU�rRs ~*�ӛ��� L�헧�W�i��a�
ڃ�VR=�
�A�j���n����yrm^�$���w����'��M� �j�B���~�4�-L�'Kk���y�x�c����s���c)�8A��9|N�[���.P
��rw~�n2��	o/�Q׺8�%`��O����8&1%�F���2�AV��x�`r#� H['���̂��K�����;�F��,=�3h��Vd��3&�ra͏j;Ga�)D����Ks8���'S�5�Q�p�&亟��򻵈.W����M�Ћ3�,@�=t���������(� ���n��&�c�ښ�r.�V��g�������)��C7������]r(Z�b��wwH��M`$�f�k:�{3N��Nm�;��k��|�K���a�E�%��{�՛��yqr�1��Bt�?0�o����5��l؞����&Fh5������O6��瓗��3��ۻ�����`��E7q�X��T�?���!�r3ݙk���������J��{y6�����&$Y��T�D����������¦��u�'��az��r���eS���Yv�.�z��G0�M,.&S����y�7�q;���c��f�.�"�)�Q2c��u§xqK�GL3 �q�@Ť�v"���]Fߑ��sGR3�
���`=��a[ԅ'��R�P�WY�U��s��aQ�I�,k6�<>�1��o�k)6��ǔ��҇a�-�O�pk_�_�Ug�E��5���עW�*�Tf��[��3W��k�-���5�
\�܃ `K�E))�q!��Cg�!R��`�LB�ȟbpW4��9y�̇��H��7.�Е��u�i��#���>�S������x�C��v��sθ��q��ɦ#�	ev����X��M�^'ƪY6��U
�w� �/�oS;���q ٗ�ě�m߿=�q0�ho��`e�4�ł�>�t���t.}3�v���"���n��'��������ޤƤI��Z���qթOA/nqn��>�|!S�f��a2`E8*���/_WӢ�*G��O�"LA�|��W�U��hV7d@��8�'�թ©��э���PcZc�ĉ��;'��B߉�����T_�&�f ��6�����aO 7N烊���ƪ<�u��t��ߙ˩/-�Џ@*�^<��3�=p���#���%��r]vH��2t��a��+���0��~�<�,�����^̗�>=��nm�:�MC"bֵ?���-Mz�k]O񣯔U^ց���.��oia�MY�f�{��N�nr
�f�9�@��5;����q�)3<���ok���rEq%��S�:�r}v��"%2�eCc�{��&������D�[�!K9n91ک�Sڐ�&���y�1����i�g'tI��m�~�XwǖG)�T��Ov�z�b3I��DN������˲�S�e��ˏ��S^ī�3�/���	�O�+���y@`��r_�t�2��P?��;!�c-���0�!��f�}l���W�y����&.�չ����+����ܠ�nO�k45צ�oi�����嘆����3_rWVc�[�7I�f0EU`���sU���Dϸo�cL߭�b�`���d�Xf��e���x���t�,ㆯ���K��9%7�*x��m�j@wA�hU7A��8I�d��d����fϒ}-��g��G�̚�#֟E|�a�+���D�m=�m�P�)�L�Y��Po���i���U�
��p7B��qp�%#Ǿ!©Q�<n�U�R��pfV�}�sX��r�Ȯ��]A��{*��z�9���(��@$�WW�BS'q.g�i��B��&^� �3bIԵ���Οx�ˁF/�� ��c�V�+ݿ�2U`���$�TJ����1n5)=wS�苸�4��B ��t�%!k�N�I�ϤA�#yc�K6�����!@�=�ݒ�w:H�YC���lkhp"�WDy��hMr-$T��c�:"�`^�uZ/�+Խ�c���ń�C�w�Լz�C�J!��/)�g;���n!�shF�����!�O�1H��53�@�S/:g���F�`�� ���>f6�>%�$��Q�;L�ĝ�۰(T�[�t����4O��x��Q*E�Z}���K��/�To�`x'�Ҿ	U���C�˛8J�e�<���0������Hb��������su��=�Tń>^�����Э������z=�򩳅2G����9��i�t��]�X��=��=��i����WP���B̲�w�wW�����M���`�C�\��Tˣ�ԩ�V��0�^�����A�R����?;��Njב�_8LEY��;�KO�\�ȍ��/����|d��)@m((��U��ei7%�A�8ą;4ha��5��)y��p�a� n|'�*':�YӇX��-�{B���=u$��Ɵ(�a�!�,y�eo���Z������CE@��c�i����s� �mo�'s�{��OYX��Q��s���FBڧ�E�1o���R�m�i�ML���x�ngHw��=c�d߄Vz20�n+T�`�;��sIs��1���S�����SqK15e')�eNK?����0W7	F��y_g��A(�Ԝ2PPT�M?����m_K��*'
Z��F�!��aT >jK�[�j����������+o�	�. I#�&������x��]4��7iKpJd�t�4('����u�[5�b/�z��⳿(M�7ͷ�J.�#MQC��&'�ᔓ������	]ه�8�<���ð�Z�X�r�[Wc:Us�6񎚌�T�� Ê�,�M�XW�n�|gď�M]�����x��}B�����]�xpgzOlr�5ۆAع�j�7����h���Vb���.��/�YV��[��bR\<�s�����FC%��/��|_?��ȒӴΎfF}/A�����p�5E�XHӎIDY�r�H ����V���k�Z/_~�#:��Ui���ـ����D�0U]4,ݰϬt��O����bu���'=�j�ꬦ;lAUw�Ss�6]�p>�� G�HF��i��kaO���ttV��U��A��Hܗ���y�	$D����#w�l��³�M����Bk+~�g-�BDKFGV���Y��k���f�>�<c���A
�99��[�.�.�
z���i�nG^o�aQ��#�`�& O0
�Ә�%���lV]�,�V��y��#�ۻ[b�q�g` �Fv�=b';��������3C����1��ZY�m�i��+GI�)_K�+-�8���'��Å�3��!����v�x.r���~�x��3d�ؒn����D����/�;��^� �]�ޞ%x���s�Q��g$NuVlYԢ �;���!��E]q�]�w��+��z?W̵�G<�V�N�TgmQ�ˀf|S�����`����������rh���=��?��������PO�lSBM�ݯ��a�g56�筡�O����������V�����q��E�\XU�Tj�{.����̙�4��s}���4JA�y1C��T���My�յDsy���ʎ��2Mg9}��^'Xi�zD����h�eΏo�45�i5�[��0�b�,��V�u4y�n�q����>cf�Ӟ""vpQ-Cd�pTv�3<{�bn\�C��ڞ�U&_埜�]A���&~�R�KK���=N�[�Ej�?U���R��܌sw{Q��FI��SkMC>&���
 �)1*���P��a����8]pFu�_�&O�୽5�í����*�K�f����C�32j�k
�̈́���3��޶9K��U)D��!n�#C��\9����
=�@�vC�W��9�5���Hy4�7i��)z���/Z4�>���eB��:�C�<�%T��%��(#�,�j<�Uό �/��E��P2wc�/Y�9t�B� ��|���mz:w�l㘇��.�����N��#�OO�}Μ␅?�TSj��ƙ��G\�E�����r���l9�O��˿���d�|�
��~��f{E��q����_�ၲ� ��`����?��{UhhQAd�E[����B�R�=)�ˬ���-��Z�#H���1';���D�H����Tڛ�A:��B�s4�n�\�|7�v���T���xuE�^�������-88@%H�<�o���u0���ȁ=O���v�@�2t3a�������;�W�,2P䨔ye�������m�+4�S3b��r��&�M�
.k8y����~g7Aj�*�ma̮YE��{�\�N���
(z�9�ǼאqߏP�qS������ԏo�{o���Elw6�:s/6v�@�%�h@C�)�{������H��/��[di�9�A=1U�S��&Gb��H��,�*�GQg��LI��`���UXR��Gdw~��� Z�E�]�N�m�l��z�S)��������k�/�3�h��	mS�+�l���1�qJ�op���?|3�!�NO�i/0�?�*@}���k"�Ԋ��N��&I���4Me�h��+,��kW=��M��u)^�`�*��՝�2��*�풢�����t_�@�����,��_�0a��mvU����?D�o�w��H)�}�P�G�30�R�eLF�x�;t�S��A�$��I���������gjێQ�sh7�� ���J�R"da�A�:n�͘-!^���{G�F�JQ�ֺ���]
�����=5[�P��DLkFջ�c��[P��*��03Ն.�PB\qkw�s��yx7�l3�<�{�-
觫X��#}���I�OrT����P]��J{��2���&.�(���$򘸓���qIkRi.ڋc��^�R�e��IςB�Q��3��a_y�����E��Z��U[h���JfĆLH>5�Z�S�Z��g�W� �C����!kg\CI�8A\��c�ð6R@��m]!;-�8�w��Y^�_� *hKEeW����-M�Ͼ�"�=T^���-+���c9[U�nz��:���;Cى�!�p3���;�=���������'�O��1cr�İ�@��/u_������3��+��x6��o�H� �;��P�(ܰ#y2���xS�u�O����h,���2�o�`�*�ZoP<'�� 	p��X�f��-s
�em|ݾ�6T���%c���t1ۜ���>Zu9��O�i�]����������K���~�p�CgWz�r;��֎GX��j���)t��3�x�z=.�W��ՈW�4��Ҙ��U���ڳ�֦�:�MR7�`�*R\���^hG�����s��ٔĖ�8,RI{��:��$@F�L�H���L��m�����Q��-	�~Fi/
��7Y�D�qm�����'�àv%s�o8��C4è����.����y��<O�n�?+*�Y�YΚ��2���6 ƑƲ�$�ˠ��$��Ģ���ej�_qO�ZyF3��8�E�Y�c�<T�.���U��;�{���Ys�Q�y}s�U�F}FC��1jw��I��(si�V�G�xd�tg���Š�=^<��t92�=nFu��&�;ح�s��	�̾��N��H�S,�v1Pq�)�� K@�KL����v	;�h((_"�gA(��P/ӄ?�A��)Z��V�E
�F�O���/K�K��>���YJ+քz	5�T{�(#���� ���\��'���7$�^e���N(|�uj�|�]0L���K�n�h|R�2��%�#�⍅F�Ø�������M�!�����!���L����m-W��Y."����ϑ_ ��H�C�KM[�O�i,�g\e����w��j`��X���]�wpb�-lͶ��A���m2��i�ӢG���Db�_�)�$/�PB�?�����\�D"ؿ�aǁ߆%T{�}?�?����:A�Ω��}�	�����ӫ�@5��H�ED��߳���L�*�#�5�~�%:?_�i�O-4�`�Yy��KP�4�b°����8��T��u���j��ۦVRRU�s�@�Id|9�� Bɪ���ͱBi�"a�ӯ���#V�x�rA����zA�{�Ry��%�����wwc�]\M�
� rB&ۈ~c�-B��K!!��N�(���D�����c��ZA%D9r�[s��.�*bꨦ���X����o�T�Q���?�`�V�Ok2��n+P%������}�V�Uc��#t��[��н^f�A'̘2�;y�.:	�"�3z0���iä�h9"� �Gׯ�)zV���.�8�&�'���P�R��vAo�1y,.�²�����g}3S�d�s�u����E�[+�V���}���7�ه	�2�1�LuKg�Ct��_���(�"=�.��]�1 �X�`w-w���eZAڵau�1�ͳm���a�_|��F�D��{�M��L8㋋���r�9�8�[?�_�R9��kKl����לB�5�Aͭ�կO�4$�]��.jr�Ѹ���~��֫�Em�X�(�T�k��6��?�a���N��J��y,�"U�Ϝ�]��6�D�����`��eЫ��)`'��z�q���[eI��������I0��P,�Z�0��y���q1�D��Yf3�l"���Q(C���SJ��&ω}�-ɸ��ɇ����:tX]<U����ER��ώ��=�`�[�%��z0�����Me.2�s2|Q�VI	�fk�׹>a������),�{�J�vH�a��E�%p!��_˽{Ʒ5����X��*[b�f��Q��3K�kXX�}�� *��9��K<=*)_��!���C�^ �@Җv 8R��D(W�8k9��K�}8�HTk�7��P��^�����7\��>ґ���Ԕ��C>	���q��}��pX�#No�����������W<��u��K0rw`�A/�T�O��,$ ��:�mՈ�g�݇��������x���*2�,�r}i�F���+��g��� �/��\^󔠣��삐b{�g��O���.�� ��|��ѷ��׺JEn�+��H�_!���ӑ��I��#�!�Uf%hL2�d���Ӊ���]8���rˇ�E�h�Z��C����'�n��������4TU���tf�} ϻ�W��7&��r��� u�%��h�#��-ӿ*@ �W<EJG����½R���䣂r�v���2�fLa�D��<����[�r�N,���o�n�+K*�7\�m�<���bL*���bMp!�k���%���G��B�����a/jpY�	�{��2N�e
í9�n,���C�O�q7� l��6o�2�ͨ:Eg���	�E:.�v�+%(`�C��{3���\����I����+[х9���1�8S���&�/���BX'�E��X�g��IIF��tZX-!�G�Oܥ!���,(�x��kN7*���y�bVSI]�-Ax��oU�a��3a!1!��	�v�+������u��,�j���aAd?7�&!�Yy��y0�}�e9}�����F�/>��	�&d�	կ)�C��+g�~��ՠ�Lg��H�
.�y�������e���=�����?_(J�������x�\�c���2��U+:�:�IoN���?���Bȭ�������e�!x�xtG���$��2p��/����������jv��
�77�
��Ðњ�"d��S��z���z-� _��qyGuZ!��!��O�W���{ۺ,=�h&P���L�&ѻVۙǾő_��/�i��B���qf	���4�P����<d�͸K|���U��}�e��~r�/��&]7O�{��{��r2�|�(�$M����Lqd�qi��݋>4^��- ��I�os�k���|-��圐��0��.��ǐUV �����J!��gB 5�S�GJ�.����� �����{k"��I	z�A�^cy[�6�Ӻ�Ph!6{~����w��Yy{����h&�jW������<-f��\";��^��SL�+�y�ctoź>�����r!�C�X�!�_G|;��~+�.ʩ�����y��;OzH�1~|�+|�@�$�/���O'��jc�`sJ�\�m6"�J};�XН�U��ͬ�|P��j�I�n�>���[�
%��%��oy_ 'L�f	�]���6d5����e��ݹ�z�IM҆��~�3�U��w�$*�u�҈J<ꄸ�(�+�'�����Y)��~]Yzs0|��G�Gx�Y�%Q��!ut�^��R�߳��=��]��TW�O���"��Sy�ڈ�z�-�u!M�ʼ`~1+\g���~��ˡ&�fô0��4P�R�y�5�`Q�ۆ����L;�-����s	����y�./e�������_u+m*����ۣ�%��8�5�4棫���]�y�n@���n�w�*]��Y�����2|���<��GR$�Lp�|q��x�b�eeԒ�gZ4��ܸ�E6�c�/l�I|,�6�5����#�{E�=Y�\|Q�GBs��F�lx�&}1eϤ#r����iڈ��$yx?��g���;�]=Y|O�:��2~#�na�V��;���s�1�g%�I˜�W-S�T�1k��)v�_K�����^�f�.		�ü�_ݮ�AC6xԒTP
�?�4�VWUs|����
���F�;�}̀�$K=\߭��D�����rC+���	P�B��#pF��[ϲ���s���7߬���`�j�T(�]�I"nu��XQy�0(�)7��?uͭ8� ��#Ól��x���d�I�CqH�<E��}F#����9	���S�h�:WG�!�Ĭ˄JN �:��~��M����d��g�&�����n��g3�3*�Pp�]*&�p]�l(�}���1܂���}驦"�b1�7�$�/PhN���U���\2�|ؚKǼ��%�ja�x"�?Fg������}%��n����5{rH��DG���1;�.+��ȫUD~ �:�$i��d������fk�4"ᳰ�('�B���-�u�ECݣ%jg(��qX�Umo�s�ӫ�xn�4� =�r�ŋ�kJi3�!aE范���V;���jA�����Z$�6�yá��.�xiwP�4��vRM����{R�B�
~&*W-�w!K�ڃ*�W�4����!��nOcZV"A@��9��
[NX�.k~�C�B����$\�o`:�Q(2���`s��O�}ʭ	ޣ%��Y�"�c�?V��4��#O��[�4���{��<���";4��U|��`-3�S(��L�c���{-[G�6�)��ۼ!P'8vw'o��"���͟ч��스.�-�t����c�3�2��0ը�:P���N�
�q-��T5(����
���og�Gr:g�f̛�
�F�1���th�i\]Cfg�S��w�>��~�uK����~���Le4m��:�\g|	�@��,>ɖx���v�f3Ͷ*�Hr��T�3.�?A�g��ن��lI��5�����5l�����;OG}5�/��I5��L�«w|��eE��X�T ߟ��ˀ���#��ݻ)���H��Jwiy'���q�W��?Di���R�M�R��2�㳽'��z�f~�&aBeĎs��o��ɋ��~0��),?�^��y�<�q�5f����fn~N"XoQ#c��&s>��1G����n^��c#���t��k�]7@C���$RdW��g�=DQ�[e%���+�!N~Hf��s휑Q5�NI�fkǂ�>���@�9)'Rǥ<+�a-7^��%�p� 6_Q)۽��5�;D׳YE*��f��o��P3�K�k�"�ͺ ���@nܔ�-K���)z��!dxC�
��gJ�1��34D�,fTWe�9������H/�a7��_���=������>�`{�[��s�CyF�[�'������ϊ#	��Ǿ��K������Ū*�p�Fsnw���/���o���8u/ j?u5�m��r�b���ywTڑo�ꄽ��*S�5Bg/�}Ȣ�{�Ќ
$��"���;;��oNJ�U%i�+�baOR9�A���|�=���/�E	��ַ_h^��[4a���~��I@��'��\urU��:hGlidQ��D+6�x?��3�g�b:Ҟ���Z4������'�Nߺ�J���TА����5����j��R_J7_��-����Pu;{7�C���Z��-ng@^n<�D1�n�>�ݺ��3pv�]"�v�vW2Ey=a��������<����lm,(�J�f����8m�m�^��bie��	M�W$k� 9�`x�/0|�>��@���hcaJ(ZY;��{`��NWs�
^�9�5��F�h����qR��8l�o
�C��Eb{�d��:�Tv-I�%�w:C�{ne����6�ڦ��U�O[�X)9��1Kq�SkF�&�B�~�|"���� gX�jI�?��
X~YG�Gn������sʶ�!eNR �br�\j-S��ȫ0��-ļ	x3J^<9�	c�+~���*/����e߇��J?�z�!􄫴_,�0s��R�}=R��󆗊���K�&�V�*����+�ˍ�����kM�+�f������W�z�֠�Ւ�͇���f_�s��=K�Л,����0�m�Uƻ��5�Lo� X¾-��ȭ�X���#E��#e��x���t�2�㷏��M2�����ۻ6D��j����7R���=�ѵ��dW,2�`�n�C//-WÞ�ᇱG�/\��2��𭔅�t������k�=k�`P�lHL!'M�י�AC�����~��d?BR#qa�k)Gk�����X<��K����!1�� �}�xE�6nr�
�5<E]���{�픳+�l\�(�_$�{�s�oq��i�M��z^2W��`OI�| �����;,��\-o���n)d`�ݐ$UQ���5�XJ�}C��\�5���SzTËi=h�T�� �i��6�k�׳I$�AR�cT�6Ȇ+�낓!1��wkr�Y�ki��kh��W�Sµ9~�-���t-."���^צ���V+e��c���U/0��"�ͤfCOG !�ܲ��H;���f�C�D�������/O5�c1��UĦP�@��/�8�����炙LI��G64�<�"�XF;�BD�^NF�#�l����z���`��n������Ƣ���� �:oԎ$'��	�ς�Nͱ?����e��ݴ�z
�L�A.��s��U��R��S5�uo�`�EG�n�J9��B��A0��4�=��s�z����;GӘ@����T�t�������=d'|��m;Wa�"�s@Q�rp���c�U�d�<:M�~�`yX@\B���x� ���\Ï�k�o��R���0�>ڂ���7����IL�_ZȜy����1-!�t�p/�Z������zTmm����`+$���%���8��(4y�7�f���'�y	|*���n-�=*���Y� ���䠯������l$v��Ww�k���xXe`�'�YZ�7l��X�E��csB��������ɟ8,�{ �zY��[Qy6s]��F��>y�1`�P��V򇞐wi)P��=^"xIeg0u�����=T��ߕ�29M�n|���;��#s�������D����&S�	�1��r)�s
KН��`���^	%�q�_��mA^m��"(P�#?Vly���0PS�i�
��%F	(���1��IKx��;G��7 ��M+L�	k��q�K#K?���������ME˔7��h����F(�����u����S�����n���"��(���C#�d߅|�E���Д�
��g��W^���Z�͂/�t��+���c��Wt���=��eW��* ��5﹁�M�dI�_P�g4�F��:�å`��'8��bw]�_�pXa^l��!۷�<�Lk[��.�X��Zb�-���/��z���,q�\����u����Ϫ%�z��s%�?���|���5"}��M�I���!��5�=HĘ�Dj�ڳyj�Ie� hX���~H�:u
ri�a��I.���1����4���`�؟=k���~gu���8�@j"w&��~�U�Xas�!���o�# 8wYO�CEiN�ha����`�V>z4&�A����0���seyޝ��b�S��w���Փ�M�t�ֶ$B���~A�-8B�K�4��e)u�����D��O�c�A[�Q9h�[)6.<����U��o��o@�QC�:��m`N!O��(����%� �}�}V����N�#*̷[��8���7��N3�;�&p�Wa3��B����^���hcGM�
)�2༜��8Q�$'?�����@L�,�M��.�t�������3��ٕ����Ì��UH��[��#����R	�O��hY�B��g5#���?% ���K\����]޺F�NpXw�%��9��u�W0����q��m"z��W�*|d�z뺊�ɱ�������A�.�el�r9H�.�0?������١�<l���n����5M���G�O��ƢӢx�d ���5�R��L>E���X�0XT{rUì���ˋ�W�?�x����1J�Xy"�X0���r�&�=D������u���8]��]w'i��zu{J�A�e?����1��y,�+0�a,��b����y��q'���`f��D"��Q�4R�d\㉳��4���ح��M�p��]2K��7]DR��&�==�a�[@E��F�����C���<�s��iQP>/I�aQk�M�>�
��ۈn)"�$� �C���aHz6�;��p�v+_�Z��W�5����Eh*��Ef�G�A3�lk�^��U�O��w!��GK��)���!�N�C}֗�g�̳T.6П��`W �9��'�s'�H
97c���qW�
������2>P���Y�N@%C�����u����&gl#�T��2���`�;�J���4��A�&wJ�/��.�c���� E�����mKj4�]���d��L�5��n����W���}���vʭ�e<^���
�6��Ѷ9 �J�Ɛ�y�ƣ��]%`O�|��k��6�|��G���/�M�E��G��F}_�̟�nn�	T3�ނ�{Kh��UPS�hBƇd��w���R���:��g��=	O��9ZϘ�����'L���u����TK�F��G��J�U��MO�7��~��0�E8u��%��m˕p^-	/�@A<�^[�)G���׾��0ԣ8��v4B'2�a�0����p���ə�tt,�ب%�ї����mwlmѾ5�Dgb��$�+��Mf��k�&q��Y��8U�Z�R��[oTaelY�,'{;o�N�_)
�tL9��סdM��R4qmN8%����oW5���^E]-t翄s:�%�vH��%�YC|>{�g{ݒb��#x��s[� �9ھz1��SF%&�)���9P�X��g�I::+�j�gX��OG`4�WJ�2ƿ�<�ߢNm���݊�7�TS�2!�c6������U3ג�W�k	�+Y���e9\�B���`����?�N"!����t0NYۋ�}زR��g������&��ե�4���Y+�Rˍ<Z����o��$\!����-��B'tN���%��s�����_޼�O����H�R�2����XUa]��0c�ou��y���P�u37��M�`�e�x���t�ё�r��h^�%�Zۖ4�Y��j��ҙ T
7��������Y|dҜ��;Zg�~�7-򥶥ܽ�G+%��{Ӱ�fM0�����0�=�P�m�L|GI��?W���ȑU���T����B�Ԫq\{����Ǫ<p��}�<Z>���,��\�?�$�}�bZ�r�a��P��]-h{r~�f�{�yi(��m$�.ƥq�7�i��)����^m	!6Z9I��I�b��d�T���`�*K�I��B��+qOUL�w����J�`�����5sTSU�l��7��e� �,�����k�E�I?��Aͅsc/�]6Z���!,w/�I�w&k�Y�{����h�m�W02X��#�-�&�ϥ"�hI^�m�+@�mc�^��?���Fl�(H�C
VZ!��.zA;rh���ߖ���{�8��O�[�1��w�!E=@w�/&�c���aܾ֧F(��6Oo���a�3Mh;8M�������x��̈́����+��d���w�FG�@~ �Oo/�H'���	�a��ɢ�$�e>�ݯ�6e�������z��u��-��`!u
ǈ@��nt����]v�ɼ����L����z�機��G.i������է%ty����=��)�=������>W�ƕ�.�#� ����j�0	L��M#Rr`t��\��ˏ�7�";�����j������R�x�+�x5��}�����L1���w I�7N�ʚ�o}./�w�h�G��S7m��;]j�Q^�%D�u8�e4�>��!"���y����ͅOnhH*�x�Y��I�C��g����O$��2���M��c�e[0���Z����E,DcNu웿x��l<���z�T�{��;YĒCQ�D�s8�rF.���1[���Z��YO�iD�e����x���gk��q�=O�*����2���n���L��;i� s5px՝" �?��Y� S]��1�U\)lc!K�|���ڜ�	�Y��yE4_SN�Ay�ZԈ\�P��?�1ҝR�KS�ghb
F~�F$j�s�]�Q�K�ܢ��x��Q�(xh+�\	��v윏#&���ѳn�-Q<��� �7U���o�`�$(�S��Οu;R#�N�Ǐ�@�.�%�ͣ��EC#9V��*���X���n�~*�r�s����c	ί�
��:^�^�
W���_���>+�@'h n2d���M,SJ�Z�gm	+�@a�Uc����q��]6��t<]`�DpS�l����r`f�g���y�3�+��<rbg�H�/���p1��G`\(}6�PE��2��%%�s�nH#?��kJ�����}#X�$2��\��5��:H��`DŁh�4�]�d՟���ԫ���~�\�:�i��E"U���3��&4>��;$�x�C�%�Cu�-����j��A���uUcbsgZ	�� o
�� 3V��?���>�ii��a;q+�aDVy�P�+cA���ߋ�여��y���j�.g�w�U��.��M�Y��1;~BW�~\g-�,/K�n������j����L����c�kAv�T9�![�.wKS�yݳ~����0o�e�Q^�/�a�`)��Otۭ?��%�d��ثH�/3VN�#�[NA���	�2� ̩c;�����m�3��H}J7�:��Ym�1�G��)����{8,y�'z��XBD����t]�b�.����j��_��3�ҕDM��������Q�8v����J�b9Zފnv�c;�=̌g���BK�@_��'P.7x��߇�]y/��Ix�w>-��������ҽq��#3���m�Y��R��|���u{���e�
vX��චO�r�f�)Je?�:�����ټ�l?��I;��M��5�N���HO�mآ�6��+�B�#�-�!�7�E>��X�d�T�%��g�������Zλ�`���TJ�`�yMf���4��Az�D_���dZ��ï��SH��'�'�Ϋz0���\�Ge�(��p��U�[�TQ0��P,��f�as)y.��q�JM��Jpf�N"��Q]��������6�����mh�A'[��I]-v����R����Aa�=:��[���+���WsK>��bsc>�Qk��Iz�(k}8�>QZ�v��)n��[��y�ac�����p��_ǫ��L�65�3K�iP+*�fjf.[���^3���k	�1��������J�!Km�@)���!Z��CX�HY�gs)X���MW�~(9 �����H�ϸ7Uշ��+<����H��F�]>#_�QL�)�sC� ���[��E���n#����AL�;��t�`���<Y�wq,�/E��HL�.f�  O��;�m�d��X[Շ/r��� ���R㻚2�K�}:sC�qㆌ�tZ����Qt��1Xc�%
H��W�at�X	�O���:��Q=|v��b"�w�E?����&_[���?�$�/����V����ӹU��mh=@dkAӺ�S��X�)g�����Zj��| �'����0�]�|�T�mЭ��. ���ӕH_�7�����1��u1�����Z��P�-��@��<V�ū��]���)���9vo-K2{��a�֌�MW�����Üc,>�� %+���t�5�m�/��xb}�h�F�oM�$Kk�l9��Z�eaF����у��a��Y1�{`8N�k
�>9�#���J�<vq�7�~1��[�	o��y֋EX�@���:_bvc�E%��CW�{�:�-r�������[P�|9�}�1A��S!
v&3W�`��?��.�g�^IU���wpX��vGP�.��M��e/�)ϕI�$N����X�	��S�u����)ȼ	;�rd�3���r	Y�+4x������ݞ��[�>�r��?hB�!*;(�U�0)���}s3����[�@U�:)�&�si� �|���+���E�	Μ�b���7��n��x�BOB���[�����_9&k
G
��̌�]<�:��㖋U���+X�o_	�4>A��'`��-J˟�>�e�8�x�XYtX�{�-�������@��q T���jG-Ù��7jS����F�dM-S���ϹE�-������G�:�6��&>؅�ţr0��k�0=�Q�P��<LׇŻ��[��V��f��J���~B��JqWg�����ev��+�<կ̸��Y���x&h}�ƺ�C�r@�
�kNZ]�$�{Me7��h^�(�(�C$^���鲿q��?i�q�ϸ^�ۈ�s�I����yW����e}t�$M�}�I���UG��뼦JRcS���5�zS0�E���9�U� ����,
kS�4IZ�XAHn�c
�76>M	�!*!'%R��u w�iYʫ��-^h�Wk0b�o�1-q��*>Q"lN^��g�+�c%�4ŋpF���ԃCń8!���Cf;Ma�ܓ��z2��������YO��1�v�ĜY�@R��/a�b� �Dט�q_���V�6jK��w���z;sw����M��"�?_����%�ߣ��l�Gۢ�Z;���o�M�'}Xq	��D����W_K5e�bhݪ���ҷ�W�3J�w�u�1�ɫ�u���;��)���I�x��7'���˾/ zD)��Z�G�Y��V����t�����d`=����^W⨪�-��;וޝ�Z��&��M�E!`o\x���Jﺩ=����e-�E�S��U�R�5Á&��Ew�8Q��$^L����R��r�^c���jzh/vs�#����r�m�ќ���Ì�%��8�-~4/;��Ԁ�
%y������n�� *.4Y�&������"7:�2��$l�(��6�����3n�eV�T�`Ze�5�-��E�'c)�T��&(�����Q{vC�Y�]3Qos�s��Fi8��h�1V�8ϵӇ.qi_��31�x�zg����>�=JY��K.�2� rn�9��x�;D=�sp?��8�q�:	��S�S��1��)�r�K�{�7��7�&	����9�_΄A�;���tP��?�?�훫FsY�
�F?����\�g�#K��ҭq����=����+�0	�?�g��#�
��<�ȳ��5���7��<Ҭ���(n�����u�K�It�A���Zڛ�H�l�둛�#tg���(��@��Z��t�����ZN��d����Ԋa�k�Y��W*��i��8G��C I�b�/��M�a��U�Ig�*����pG��V>3�Ĵ$���]�2$pN�l9(j�-8���餱~s|�����y�b�Q��q/an3�+���b��\�z��+�;�m@�%���i�j?W�5�&8��`�}�k.����ӗ#q5LBH���D OV��;�e6�o=���d~���:�5i������Eȹ��|l4�Ѱ�럳K��8u�т�Vj�t��*'Uދ�sB���5u}�ǥ .�3����X�i��a���<HV�XA\�cA����f��g�y����)�	Yw�`�ɋM�^���Bڨ~w?�-.7K�Ș��3��[����L�}�c�&QA���9^o.[�v.�����y0v�5��o���Qy���[`V�OW�ڵ�%����3�s� �V46�F#�a�[��ֽn�/�-+����;e=/�����3���k�ե��Ti��?TGÊ)�a��th8*n'�s�������-���.��L����:"3?X������Z�ˣG5����^=@���Pؚ����8)�g��~�Ҙ[�,����*K�u�]���D��w�TNʯ���)��Mk�ӝ�$���mXYF�M��|Z��0������n������RroѶ�$v?R���>��O�l�S��$�O׈�25=���9�OXj�I�ޚV���2f�6���P�E�X�RT1���"(���әM4���i)���+JH�y�~��ψ���\{D���?˯��njׅ��'�Zz���w�fe5}$�{�=��2b��0���,P@k�S�yIbLq��T�f�l")�Q�!�7�ۧ�����X�b"S�|w���](����CR�؊�\�=��c[��i�f����5v9�w�Hs�FQ�N�I�x�kXC�>M�r���)O�Ƕ�4�a~`��1y�p���_���h�5�����{�*G�2fIɉ=��3y1kD7�͋˭��E<ܥ&�K(&)�4p!�'�C3�O���q�$���=�W�+�9J��i�H��L7�g0�����M��>>�%��^���C*�H�,/ڸ������#:�s�t���D�S��8���s��7��w�.�/ b��Mۤ� �S&�m�@�SɊ���]��;���d�����
m}����l\����Sy��lO�Ѭ��� ��!W��d2�SdOccor)��l�|�yJ�=ې��K�E�oD���_y	��A��?�t�g�1����U���h8��dbD��u�8�ɳݩ������T�Z��weD'�Z����!
TApЈ��i};n��C�7p#��^�6�L	u�;��\x�Q�-?@�<��o��rS�.rK�������v�8�2q!a��4���Q�m�Ǚ��:,��l������u���m��xo�
b8<0�a�.M\��kґ�| �O��sO���"a�"Y��F{�p�N��
/�g9�JD�WQW���{q�@p�]M�6@�o�O���ES�i�u�!:�/v~�%~�C2��{����� ��}�fZ�[�,9]L1�XS��&n���OU{˯��g�ѦIp���`�%X�T�G��\�����T���e��N�>9��F�A�S5�5���jȷ'���A13M�>���	�D�+������x�h�Vlh�͢�?#V.!E�r�З�0��Q^�}�;����K����^&��.՛,��k�+S;�rQi���h�<�p��m�е��+�*Vi�Q$i��ф��_����?�! ��H-�w���1�U� ��&m=o��d��}��_��kH��z�y�VeS��x�8�t�p�����8���u�L�����j��k����7ct�nZQ�T�d�ݕ��H�� E-(�n�҉�G�oM��t��A6օC��M�Lۦ^=<��P�ϰL2���B��3��KK��w`;�Ux|B#�qRs<:�T� 
 ����<PAϸt����ee�˛}��O��r�D1��Q]#W{(����O-�8(��,$�������q�_�i��%���U^���l�uI�c����ڢ���_��)��_��%�a�nUB@|�F�}J���j95�KS;O��p�%e	 ��G�dk��IuN�A�v�c��a6y`v�9!"�P���w��SY��D�w��h���W�N�
�s-
(υ��"'��^(����+�p�c`��&���������C�Ӻ!"�-�;(zȺ��
���M�Of�1ꇓ���@-t/�6���Ғ��̘��H�.6�G���@��
};��X�/��
�}v��N!�����Zn�s�q漜��vW��O�o���'8�g	��ۜ��-Ј���etʯݥr�s��r�������1�u@��6��$�?�{�ѓ�7ɲ�f��Ժ�jv�z�f0��K"G�i�� ����tox��z��ߟ�=5�g��A�Wr\��Դ�V�F������*�a��MYY`j��\�]��!�X�ϡ�� �� �PRP�e�!G�ֳ��i�(xL'�h�-np��<c�}T�e�/�/k��2��˱cm
���� '�ǘE%z]r8��4��죗�o�%F�yzd񛃟�nޘ`*��jY�٪�����ݔ��M�m$�n���nÏ�T�ΘjeQ�8BsZ ���H��E"+�c;-�5���Gg�D%I�{1�JY�H+Q���s� F�Jid1Q����3��,�izr����&x�C�g���ŧ��=E8�ߦ�62j��n��B]6;��s�.<�ӯ;�5���=TS���1׍g)b��Ka��r��� �	�#��/N�_�mA��]�~1�Pv��?���HMA�0���
���FZN|�i"�B�K)�6�.������,�+}�G	����{#�i�G�^�c6/��V+�7�����V;�(I�C5��uqk�D��ic����Q͙h�l�#����MZ=�嬽��lj/��=��iL
�^���%:S�����T��W���J(�0Q��6�� $�1�j�KMb�T�P� g#l��w����K2���`ß+�<��]��{pIh�l����/ƹ����E����xb�ۊ�X�/������}��\�����Ǩ��%[if�d�m?�f���E'�0%}�Л�u�ҖO5��H��D{<���������"��| P~�8):F{Gi���2#� �á��4��M����[0Eu��%I�QjS#e�ݰ UY��s, �p	@@� )T�j�m�t�i���a1z��l�V����A�@$�A 6�"b0y/R��U��� w<��d}�M�����1B�);~���-�amKhB���E堷|�����`l�cF�A��R30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���<H����\F� 8�,]�(��afR)�a�sv^\�!E�׶W��ڮ�-```��t�q�8��^C��YuC|j��?�9 E~�:`r�Ķ12~Up�{��Z�z�H�	$v�J3~�qY]n��FuY�� ��.�?��7����
|���8!�-��F���+%^�X&I�wWB ���A�����
�t�-�ҤP��m�͖���x��'�Ŷ|�2�93��K�����fb�m[&�2�Nj?�Nz>��9G�:O�j�>���G_(:�^E�gT�u��G���L 9I���6؞�|!���;�tT��6����9���ܭ9���E���!�'fk��3�rw2�a�W���O��x�����n�ߡ��H��g����-�HM9��·�%�W��Y?_�-#�'��N�����b�!�Cǹ���i����l�#Ӧ0Z����.0y�b��9��mmtM�ŀ�n�o�(�i�]ȴ��I��@�cw��:J&߂�;
a#�IN�CO-���\s6w�;�	+��=��[S7a�$��c���dJ]��}����(��nG\\�p `/jcL�����D���t��<=x�~e؅p.\l��>�NE�at���;Xk����=���q��,8���ң���z��Q5/�����ė{�5$.�E���@�}��i|�2�o������/5$��ɷ�Ѷ'ѕ	�k~w���I�z��6������B�����̀�I~�'�c&{ƐN\���Rؗ[}yu+1�=�P����{�	�:��ki�w8�؍���K��j'���z62,P�
^���Jjk؞w4@v)g��rz �!�2�� ���3Dfw�e�ٌ]���8�@�d�S������܁Y���KG�ǧ1��O����#G��GB�BY����2Qv+���.P3~&,4'S��&/�q��;�a!�@>��Ik�3�K������D�'�VHN��@]&JeO��pV71����R=m{�D�L���?��`A��R����#hD������@b����NK�����yL~��Y]��e�93?ix ��J`����P�N��05/���e�	�N�n鯪���@U�K�Q)��',�gK��=yN
4�3W�`��.+�t��V�I��w�pה �"(�ƙ�
��u�����䨜3��4+:*�Q�ת�,��	�u޵�:��2G�RF�"Ofd8�NM��"gI�kҤ��z�\�o}z'mO�=TP�硶�����o)H6�/M�\Fj��9�͔/_�iH���)�yNn��0�z�4����Ć{�]���
�f1����D��B5�T���G�Ump����P>FOeL�5ѬעSm�.�vj)�*K9���{�p��$����J�f�wǶ8Q�j������||W����Eċ����ط���vX�	��HQV��'�RJ{�ĭ[�ii.{V�!�5�4E���4đTEv��L7c�����>k���l�Gs!�H��0��O��
xէ2g��kcc���, ����|�w�Ev���!�?xk�g���W
�*i�\�Ҽ!��9��E��f
��=�_�[*B��]��w��s7�-��L	��O-,{�M�c/FSG$*qa3�!W��a����j,����-0}�C\�!����������>\:��?��J�K��B�� �҆Ts]k�:�Q�Q��\��| �����ӄ��X"q%ɻ��S	��Z��c����{nZX6r����*�.:�h����
�rߧn)�	~�㸇ꁫ$:�ӟS.L�پ�a��ږ��=�(#������Wb��a�T�"�M��~�9b�
&�']��K%0O�+=aO�>�3o����';m-�<�7�������ɍ o/��(H�N��}�;����9�Tw6LL6{&�VE�H�^�mF���o*79�L��3��������y���=��l�K�p��ʢSJ�󃴇��S��P��B���hw�HSA$���YHɝ�)�92f���W�^N�6E�mn�^Vw��D���_[����T}H����)�=�TV;y$�h��8���ɰ��Qtr��8�(��O�����}��ʾ8i&�iբQ�BY�ȡ�T
�����)}QA�B���Oh�2N��W�ت��
o�o����a�քd�E9��_jW"��\p���z�2[11��2�>�d�w�	�2��3R�<���M�_1
}vS��ςDx9�>����ģi�?��]���KY�X
������	]�6��c�kZ�&��I�=o�����	nzfrj�S���� ��c�/
���$��^ܱ@��rZ��׫'��C�#9�7̘����ݿK����5���PÈݙh�dZ^�B��q��b^��{={Ep&O���:����ޅ��k�-�Es	v�t��&��sʻ�8g[[W��<�zY�!��ysj����Ŗzz�ա?M�
�ͷR��(ե��r|ԋqd8|�-kٻ�-M\^ �$g�{��b'H����_��?��w�y=��b4�
�U���'�	6,���y�;��Ágv�-�L�4JFgٓlH�j%�)������b �/8F(}6ӌH�R�.��r&ܰQ����s�8�Dr�>�S�Q���q�ۻ�7`:>%-�+��|n��4�?"��W�2Xi�z��:���Ba��#l�;�	�zC��� <�E�5�1��F�/B!hX�L�]T=��M��G厽�s�������0 4�i�Ҽ*C�_���|A��.\h�HHT��w�W�*i�ܮ�:ׂ;�䣺�V�CLX7D��*����� h�B.'9ilP������C}2��(ߵ���7T�����^"�]P��Eut-��^A�"<����|�r'a����%k��I���Sfx)9����E3��B��[ �G�%
�k�g��i��Ia�V?��> ��w��J�̜���\zu��;^�	��΢�ѿs��H;���j"�21���-�-{�^�W�C��IpOlF��ʉ�PE�YJLʫ�L?0�?!��V�Np�a�F�t�%�&�� ��JxK���S��1΅��JH\�W�'V�U~_�3�2	���w��G$�	�"��l����f^�_Q�|d�I	����dq�9>Ħ�稇l =�:����u��ȟƫ	o'�X9��~�q��͖��a�O��'�Ư�����!�|�&�}Sn x��^u�P���U�yed�$W���vB�.7�\ 6,&E��6,��(z�D[�4)�I{���ܿ��>�����5%tH�(z�Q߅Y����r+��>ԕ���2��Ǫs���<|X%؍�bb���d+y�Z�f��aEC�.�F��P���f��:s�Z_�^��{x6�|jb�.�&�<^K@L}_ȣ��C)��{a�# ����o����y=U��iv&��� �in0�ay�u�T��MCU$O'��&�B%/ȣ��'%���G�U���5����N<��]o�/t��4�o����S�U*<	I���La�<�+�鞃΁���!�疒Ѷ��`�	���N�i��̺Zk:�����0ͥ�f�{<��'B�ǂ[W���ב?��C]hB�5����=���9��d�+F@��do��Z0�J�a�+���3��t���-#�����h��^�LJ:���m�\�D��)�����`������E�c��2��(�(q�,�2�(���I~�l6���p1���'_Pl+qumĶ&yJCY�_��#�K�hLg��ik��5��	/��X����;��K����`���M�\ݫ%W��f��X�;}�%��=�Ia�����^%J�L����*d]���)�M�LD
��D~�@?��|�c���F-8..�Vl:TQ�v���X�q��������4h~}.C�f9Ͽ�H��z�/ٿ&�X��*��ֳ�!����f�I�K��xx�Z[�G�<�uТa<�55�8�8�2}������,�Π���ӆ	�N�2R��P��S�	�<���̍R��?_��^���g[誡�!N�Go�,�~�^%Lts����B�gp�l���������A�����tEڶ��6���\ +�4Re/��A�"B���~�� �0�~]g$j[��%���:q��^�Q/�(�?�T��V��5*m�7,.��ql6�A�(�
M{�`�@ <��5����c/oK�4��֯v�	�ƨ�����Py^R�����O�����3!�܂}7���/��YL�6��!m�`w%����ajV���<�
�ۑTn��M�<�6�������՛��s�{�j��T!��"���m6�S�޿H�؁g��2���a1	t��Hl\R��8Ī��y]'=s��>�v��A"j�8�5����I˿�]�e "!}/�G{.-Z7<r������0O�^F�-^؛S�YD)oe-�\7��<]���`����p����pP�D����/�>ֈ��	9��{�3���+�TV� ���XWb9L����젊���U���m?��M�϶����>�-u�����p:.z=����l��L-��3���#C$����e�ڜ�Rs^�3�����8O�۱.��˖!]���'� fv�RC���_�d#|���3���	5 �\MR��U���:�0�gy�%:�<ެ{S�Q��>�D>��|�k�g�Ay��2���K�K_�喾SڙgT2c���n�����7&O`s
�9TS�؈iܥ��/dZ��-�*n
��`q8'����>�Q�>�v|�0h�-]�������X��M��$鈄�.�	<s̈�k)3Qpn5V�D69��jY������6���æ��(�ަ����vOn�d�ϲQ��%�q&�@��僸2�>�����h�n���S�����;��1*Ȋ�Fi�a!��y@G���S��R����ּ���pr���Z�����z>"���Rk�JZ��g,;fZ�o�Ҽ��_"��|�ѓ4^4~ӊ��| L�-UoF&tps���� �גI���
`lJ|zo�!ͻ)�['�ԩ�֭
t7K��I����7����Y���#��N$$�*��*���߭�R0��0nQ�:��#����u~2u�sH4����\�9>��0�q�U�
��o�~!�0Ɗ�pbka���Jª�"�^�HΞ��׳�^X�A�U���	N���;}���_�Y?֛�8B�V})�j�h��)�!�1r:�s�M��^�vnaqU�c>I�U�S$��%��>˃�D�����&Cc���>E�#�\{PP!�o�ǘ	>�9\��W����D���ReBL�q1q���½�*ɨ��T��� ���!��euCo*%P7&6S3�?�Í��N�NW�5Y���1�L�m�r#?bE�D�N^��J��Iu-�D�ڄ9L9��eeJ�8]��z�Tߓ�&fwH^,�O�j��E�)�� �Y�8a��P��������AN q��sn�� ��x"�1E��)�)�͗�t[� A'%������JK�Z���;R��Ͳ�y����]���w�s��F�(^x�Z<�3�ʿ�l~������.@��碶��v��s�}�DH�8J%�����B?�:�@��YZo5F��%�uO�Mo�d��[r���eS�����[���\�^����� � �c�?e��hH>j	8d�[Rb2�	w�dl��`5]TNv�<!h�Pt�������Y��������%5`��ij��sh��L�����W=�'SEv�s���q�=d�J��aH��@��I~e�i����������ԍ��v��}�~C����.�뭻b�1: /��b9�ĝvo�H[a�R���k�_�ZЏ��qlݮ��H��n��Լ���F5��u���������bu@l��#j*���o$�}��b4�o�3nXwY��j�r*�l��Kfa<VTۦ�T���ȥP=�w~^]|P�ɻ��g�Q7��n��Z)��T��<�P�S7?�*Q�䗖cԌ#2���A+��r,v�޲�������%8G���z�+E3���j}�<�<U�8�F��8��b]GQ�ʎ�g)ΆђΆ�s����T�n��ףw�ք@��Zw�`����)����'��?�C�$�,�z����gT�f>1�19p�9չ��Rz����ů���~%C�];|aF�)g��T�ۛ�Ut$�q%y
	��e�^��AFf��+2�}X�Ew���n��A%�L����~���]U�mM'��mx�����C�2�f�����Q��swhmݢ2��?�d�>i�G�J�7֢�I)_��Ctr��[�-Tg�uy��G��+L����ثW�!bs��<"T�D���96�f��ũ�����.~!�|of�kW� 	r����\��PK��,�����p����@�������*��e|M�K�֔.��U�m�,�C-�������[zbE��C�<#�uN��3zx��M������9j0F̹b%��ԭ�tɎ�^<Լ[�1ݵx��d���Rk�՛@�`�����JsS˼�8aa���Nq]-�h�ɟ�w�� ��&kΊZ�[@ҙڱ�Ic(�]d�#����V(~&�G���pF��d�cyo�註��!W�t��=�-~�C�p1O���-{	�aAaʨ�X���|=S�=�`�ڞ��N��DM��A��p��/�|(܎4�{К:$dEb��ľJ��i飋�|�u�L�
�͑l$�B*�D�j�9���֝�~�~�V�w�K:�6����� �B.��1n�M�9~ �c3`����/�� �؄AMy���j&�P�P@��f��-O{�đ��zA����+jT�k�GnW2|]�i����j�.�w!,�v��k�A� ��2,$����D�-�PC�J���~��mzۄ %Cь�m���Yj��������1I���dX�����oKGO}YQWK���+ϔH��3���4�~����į��lnnޱ@l����|F3̎A�U�k�h��D�7sZ�NG��@JWne��1ҝv+1����{�6^�#�"����.��Zޅ���h+�W��M��i�'K������k�7�f�r9�X�xA*���H��b�;Ι�:��̸veæ�Nk���������3)�>�wjE���Ȝ
/�Nw��3dӇ`FfHx˨ØI=��H
 T�K�3
��% uH���9a�������:W������s���Du�R�:� �G G�Fo�O������V�1^gV��|��B�\��$}^�O��T�'�#���7�)�]�|y�\3 ���R�=i�a���,0�$>)�-.n4@��m:zC��������̛$.`�,��%�4���"L������rUo����Y���i���9�5^�>������Rj�ӆKF�i�(�ɢGE���{��� �8��j�L)��IK|�z��E�x���s�T�	6�CT�	FH^:|�b��R��Ě�5i��V5n5p��������'��6dZcmm��k���l�=��eNUt0Q%HOݣ�x�E��Z�k�0��3��m|�њE#3ˆn�9xX���j�
�Qi�L�)"�F�kE6�
�&�7����&#~���J�y��7�*��^0���,h��MPv$s��$��qz�4�.�:�?n�!�8,r��Ѻ�p�������C(� 9�Ʃ�>�?��,[$J,�%��`���ۂ���	k�E<��*��7_f�il��Vӱ�X�Ѡ%66��`���#���z��d�^�r#b���z�:- d�b쭳0�r,�"P=~L']�7��v�:e���3L_]l��m�ǹ���O��L���`��M��o�@a�53"D���>9�r�&2�jݱ?�O��a�U���r�3\ꖲH
�;�y<�	9�d���C5 ʣ�H�H�錵v;C�x�������LYl��aVc2�H��^m�6ڜ0�9����R�����q�������m� ���x��py�s��nأ��4E�S1�����)Y�o�ޖ�VkA�����h�J�W��V�p^D���Ȏc�m;V�(�Q
Cɡ��ޜ���^�������
g�Vx�;�h�� �<̊�z�Q�D��(�Ԋ������B�}3��DS�VL��/4�B�ൡ���
�����O�}��(BѠ9OU�3Ne�%WJ��w��
�Io�qz�q�#Zd�Ŀ����WO�\=�t�D9��?6M1x$��`d��$	�c���a�	��[�Z(x1���v�^�YH��N�=O���������v?�ЦT���P �>���Q��z��](�O�����1&�o6�=�k.���	;"zr׏�S��.��S7�K*��%��N���@��frǝo׸�[�/Q�#�K̅���!���x�ē��h�4P��H�29Z��g�/~�q,�5^�=Hd#&�f���0�<�x��W�k�x��=^�s6L�t�/-&���~�8�WW��g]h!:g|s��4������F��!�Mn���oE����8W��d�q1�cښ����j3M	=�6;LTș>�H'=�3�Ĺ��ri5?����T���X4l4���U.��'T�,Z3�y����8v#y�e��47�� ��ƗLH���ǎY���'2%NFu(�y]6R�w۟*J�}ۗ�R¾s�i����B��7�>O������`E�-O��j�3������D0��Yz�xRٗiB���#yy;���z�s������_��^���B���Y1*T�6�|�4n齪��>=��^���VO A�i���*�*����A�Ɗ.���CW���W��i� ���p�;٧ĺfw�Cy��D�6.�%~ ��(?�'���P���2D�C�A&����
y�T�n�imP^owfPt�`u�t���An�ǪqH�����ԛ�Zso�$��{��@x�L���R	D��Y�[Mll4�%�����i��6�lIrF҈!�э3��*����Y�n���u���^MQ���z�l�
Е���"#�J��y���^iw*C��qp�p��N�=S�Y��ۉ�0T"�5�^�[Φ��V��7�nFݍ�J�ed���f���	���aQ�J��%W�S�VK�_�*�����w��$e��o�l������-_~vdM���U3�qrs9���4!�l�����S�ݡ�B��l'Z9��~���젊O^4|N��zh�N���n�)ly��� e����}J�"Ђe���$d)x�#|S.�]� #�bE����.~�k�zL�[�)��^�C�?I������/^��bJ�H��#z���ߒ��J��+4Ԃh�������������dX2Gr��S�b�'�Դ�tyR��f���E�.TuO��|F�g�A�^Uks�'����{��J|7��.@�IG>@�V�_����)p�"{�N� a}��O{��[U�A����E���+��R�(��y�����	��Z��U��sZ_�'�p�&�d�/D������[m�G�u[��W�� <�F]�}|/��74ʥ&�l���bh	�?ʙ�*<�߬�v:Aή�.��yz��ݟ����	��NN1� ۶G�Z�=�>�����p���{I�6��z��ϩ��
k�d����h�.5X2���Q
���*�X!����Ӓ邑��'Z�J_Ż++�<��
��;��y�HN��=�+M�J�i䯓�i\e�o�v�פ�ʬŨyN��%I�0>f�*�(S�q�ٯ2�j���@LI��6��(=�����_]t_q"wy�s��CF�}�tj�KHߴL4%Y��B����Rx�/�V4X{\���HIKٝ�-VQ�CBB\_ %i�fk�7X�*`}�]�j��I.�p�2]�kA	%��\����d��|�z�VQ��ٺ�bsA�<hĚ�5cY"k���-�h`����f�QCM���b��2������V)��L�aѣ}�ѓf�7��U�s�'+&��E��*a�>��g�ڼ�fJϟK��x?��n�bDa�-k�bX�8���>���w��
K��´���x���R��Ǳ�Y3v�t�����RI�_Ͻ�^!L�g��[�w$��*sT��,@*�˫Fmt`B�Q�|g��ElM���V�����AN�T���t2���e+c<^�)��Ρh�/�ٚA��!�H�J�Hp��3��ѫ�c.�-Y&���������G�(�a�����4)�����mjj�,�k�6�6�V"( ��MG��mN5��T�)(�c<����H�#�T��,��5���)�8PF�Z�)/��\qޔU�r3nA�ov7�M�.�&B.���!ڊ�`��8�K1&j����)#��h�nԸ�Mȧ#6�n��P��/|��|�{�>��千� �w�@6������Hj�/g˞��TN1�A!�u�t)�
ե�'���]Ԋ)�BBc�������"�O����L��̟]�"n}F/�Q�.�W�7;u=��y��4!�Oդ���eƛ��D���e�*�7 ��<*z������s��ҽJ�D��鼨pֵ�K�֑>�����ެ�ؿ�V���9(b�J����$�m`ƞD彃��r��l�������ꙺ�J�&?�p�L=QȢ�ަq���|%��>��uʊ0R��l?R�'3̀pŌ��(�&������P���( 3�BR��Ʒ��dб�C�����u͖'<�����w�0>!0�ؾy�p:H%{�hEQ�Ol>f�U��4�tg�oy���Oj�K��.�r�S�VT��1x'��{sU	7^E``:�O�KSH���U�d�l�dg]9-�0;nW��`^	�-�!�9�Qޑ����5�=��-
���R���;��q��x�QL���M�^o�5G!kU�>s�5�7mc�?�t-Y4����^����B���F�y����C�7n�2�Ͽ�����&2R���Z2��(������n�S�':�r?E�(c�wm�iSyϻ��@�%�[��_�畔���	Q4�]���rZ��ӹ�&�"W@%L��?�Z�|g�?�f�o�l�ߴ"��)��#[4ƅ��[�|�����o���t=��Ggg �$�I���
�0�|g��!Z�*��I�����*7XǃIx)(���%r����i#��}$�nE�.��������ccv0����@#��m�B�"u�)<4�<7�	��>,ڜ0͖cUv���n!�ʸ�:D�kn(��T�	���7�Kz��+�����Xޜc�¯�Q�P�7;�l��L,k���e�&�#��)�w7h�K�����r����I�n�v�$Upt>�(`�`�m���L�F�؃�ݼb΋S�p����>�^#��P��lo́��s�9�OȋL��᢭�^%(����e�ͦ�څ���l�B<�*���!{���.w^e"�X*r�k7��6�/?"���L�>���>W�� F�,�{L���mhi?�A�Dzи���V�/l�����3L&����L$ެt��l������R^y^�� T j����Lߋ��%��V@�]�C�j�z�'�G ^�� �R�-G�x��E:���d�D����Q ���%^,��T~���ZQ
m;_��_T�\=�JI���ӓ�(+k�Z�G��יl+�~�4Դ�0�t�X�(���@#����8W���ymLB�y�-"]Y���F.��%]b=�Ao����HG��(S���`b�[��-\d��	L5�-*� H��?�3Kh5Ї	�3�[#��m�x��$]l��w5
�>v3�#h�Ǎ+ԯ��pY~S�閣�v|5�6���������uŐy�|��7:'`�y��_qsA,��N=�22��wE�a���E���$#�� �����K୮0�{�v({�@��m��..eJ�O1]:�/yÏKu�j'v��5[nꈕ+�r��|�rq���@�'H\vAh���D��?5�������G=�b�=�TuT*(F�h�*�bb�c�o	�in�w�)��7��*P��Xb<��k��Z[��ߜ��1Aw��|���(���:Q�UlQo����) ?+�IY�	N�ރ5�?�B�QC���;V#��i��+��@,�e��H��V�R�9�84�1ٝ%j+rPڰ��}lYz<b[;��|Fh#8�k�]�9�ʻ�)��˒;�s�${�-ʻAiא�W�f�߇N�`f|V�K�Q���y�;�|Ca���Q:J�ߔ��3x1��p�]�A��z[���'?�d�~R�r]3CFO��a�������n�^$
��H��=/��LF�\4+?T�X��w�&�[+�A��'��Q�`����jm�m�@��*�U���8��iL2Eʟ�Q�����ۀL	m�S^2f'!?�:>�_	G�������@_��;!Fs���QT��cuv�G�L��/�_�ظ�E!���Ղ�T�T��G��P;�v7��LX�:j!>
�f�v��r2L������m�������h��K�;�1�C�6%��$C���.MĴ�����]��m�-=m��>;��ww�b��uC�/�"�J������j��J���l�0eab�~����tv���s�H��BUԯ�t���h�#��@�ωL�J������a=0�NE^1-U��6�w�o"�c��׋[--��>�ccU��d伍��p��>�(+?�G��Np�=+Z�c�K�uH���}5t�[=u��~�n�p�Ǖ����a�����^H= ��m�����,�b��ȿ��Q�/��f�;d
{��$�:E����tiV!ڨ� ���W���$��#��ܑ�f����}~Q��c����#b6 �ü)EB�5`�^=���~��c@␨�� y�q�ry�2�˗�	P��AzdA�#����2����g���enCj�aw�f�2�N��n�MkjE�wvvCb���/ �K22�2����Dqa��c��7
���V��W��M����N�YH�姠���1�����`�aA��ܓJG\l�Y�n~�̫D+�K����3ز�4�j� : � �������r@Y&��cNs3���".��?D���+oN��\@7H(e"�)��V%1�F�,��{��|�;�o���ż���)6���hލ�����Z6��(�KR������g����3eL92�xH���q:���(�ܙJ q��/We��N؛��s%�sc��.�+30m���3��N�+��[Z�w�Vn�V��i���*Ө@����l�����e:������n���J��ZU*����"�.�hh����Zޏ�g��f�o`Ћ�P9"�� ���4��k�ȰY|�e��P,o���t�~��z� W��Ir�
��h|x1�!���K����֫�N7	n*II���u����L�v#v$b��ֿْ��n���lzT�=0l���J�#,!�����u�@q4y%����>�0ލsU�����X!���[k2�%����*�\�N�\��1��XOgT�S���/��!O*;���]%�-.׶dܔX)��Uhw�}���rx���ã���v�NmU� �>GC�	t�^� �7K-��؜I�����;� �>Cz�#��P�;�o�����9�M����{R����A(�QT�e�G���/���Z�sۧ*Gpi��M�&���F:e�*c5z7$�6��?s)p���}��_Wp�P�)���L��m��(?�HtD�����%t��n=���~L7m�#���٦����R���?O�b^j��Uvj�˶�hf�>�;�6x��)�;�+�� o	$�1���~��x`�E���������W� �k%��ܒ`;�6Z�-�;G��0��M��[���5���$`�(���Z:l���P�l��6�[}�, �եb�y.���Z��B�N8���J;hB}x�>��YF��%�z����or�v��Vx��{S��ґK�[��\����s���CK �y?�},hFX�	���[������߭M�lR��5�t�v$mdḧ�\���ImY������ҧ5ޟ����y4ʈ�F�"��-��Ub5'
�ԑr�s2����="�������maFF�x����x�����:��|�]�p���F�v�J����d�>O0.�2�`>K:��(�����Yvm�[�O�f��+Ѝ|aq*k�ÑG�H͖3Җl�zEu���������x.qb�#]��vw*�u<��ӝ�8pbr�oo�,nΡ3w�~���F*�EE�	_�<�fx������2�e�w�}�|��ɹY>�Q�/)B�W��bs)Q�ң��z�*�h_?��TQ1���7#0��%�+*��,RA�ް�]�ϕ�#v+8E���;�+�,��+"D}���<"���pFY>�8���]��8*)����sA��sʬ��ס5.�B�j�ج�`פ��ܶ��q
CZ��*��kC���'V䤁1��Ip�D�� :zL_�������*~��3]y F����˫@�Y�������o=$
ǿ!���/�84Fd��+�-XQ�w�B��l�<A��ݓdC��$��k��[m�c��:株�����2���t��O3+�1��m��2W�?���>'~�GJi��u�&�GU0_J[3��d��xT
�Qu75�G?S�L+N��C��i�5!�����"�T����I����Y��g���tK�!1xf��v��rcM�� #��~���Ǫ������D�,>X*6�g��u+��8��M�+�m�PFNm�*��-n�������J�bCΧC������q؇� I�{��+��0��b#�ǒB)tG�����Y2��s�H����!�{���@��t�m�J�m���4anV�N�J�-�q0��w�F��4�����5[>R��on�c�b�dU����6�(�,eG砀p�j\��c�����\�Ĳt|�=F�z~�w�p�J���1a0�ʦf��b�=�O��*�xO@h�}����n��/KEb�q{�	$E �;B����i�jШ:�S��I���N$�XV�����۰~�c��=���V
6�M��T�B���˯Ft̋y~"�c��ܐyG;�؂�1y�`l���#PJ����ԦU��������x����=�j��ɅŽ2z�L���%j���w��vtґ>G� ��2*���s�DB���t�H9ͭ<�|�@�^8<ъj�K�,Y返�5���1�uI����CZ�m�xGϝY�'���~�+�|�����3)lO42NE摋��Zd�f۵��@jؠ�B�3Jx���q�fkvD����f�N��z@H{�eSA ���1�����{Sd�e��`~I��p?�`��o��hO��U��H���KCV���D%�>�������9��3x�O�uo:����9�ә{x>�J��eL�Ni�~�u�e�D�D�Gѓ<j�5�C�s��H2�Nu�23"��`Ĉ��uj��R�I���z� ���1�?��ͧuƮw�w�u���]��:��L��}\q`��s�u	�:;/�G�<�F-��O���'��Rg2�������\���}���O��\T[0�!b��z�)s���cd\1R`����C͟�2��-[NE�)*fnr�����z5�l�C��˶��o��,gȑ��0�������P]�E� b�Um��~���{ ڌ�7�O5�;��l~9��j�.�K^bݦ�٢�����_��eͷ"BP8\�`j�Ũό�|�Z�8��v�C�1x��������	�5H�^���
RճrĘ��i���V��~5����6t�i���t�ck��=�Qk5�ZlŨ��8���0ϯ�O~^x�g���k����h���!|���E�[?��,3xV9ĝ(�C
��i�s9�'>��	E��l
@����2����4�
j��w"�7u�1�w�1���,f�Mr��*�$�qx�ڰ쒪��Ӻ_K>,p.3�xY���,aN�����N��DJ>����*�J�L��nm�+{��W2k��u�|i�um��gB��F��/�QX-χ%4�G���6 ���c���Xr�ҵr�M6�5�u:+�u��1�rjnqbe~
y����L)0�:c���͕�L�u���
��� �ZF���A�xv�K�-��a�"Z�	���n9��8&��'\�0�Ow��az����V33ZVd��d;��<��b���ݛ ���@$H�E�J;��C��4�����L�<��V��JH��m�����99ܧ颞��UZ����(�����]��9�p�ե�������fSo����7@:�����Y]A��΀����L�����n`��Qˡ��[�my�BV�an��B�������~]�2��1���Hn�Vv��;D�dh'IƇzB���Q���D�(:�������)}�>���T����B4���
�͎��p}|��BӤOS[N#�&W��ص��
��#o�6��6�a�d�\r�CT�W�S�\{*?�B����|�1�B��jd�I�	fٷ��,y�G��}�|M!15gvvު;	-w�������Ψ��%�4B��$���$h�����O#4����~�]&|�X��喦4&V��48=�{3�]i	yr�nSf���I�񪉐'��߶ןN�	��@$?rŚl�vP�����#�Õ.��[���N��ъNf�P�L���Z��E�-�/q�J%^�Δ=�u�&�L	��:;����؆k� (���s��0t%�R&�����	8��W?5N�e�!��Ss���Ƣ�"���6M�0�X��������' �qo�KژM���]�M��jtճR�����'�ϨC��p?�Ũ�ҝ���,�4���U���'�K�,�~y�����o��B£P�45�@�޿T�ⲥ4���F��xcK�I�F��D�w��R؜��^�ܻ~�P��se�ڠo����I��<���-?�f\P`EFT-M5��X���DL��7��B����z`����B�	�#7�е4z�A���Z���$�܍�Q��B��k�6�Th�����2"ڽh�&���*��y����U ��i�:*δ����AC�p.RS���l�W�g�iل��X;ח�$g�C�q�D�l�#=ۥ>9�9''�E�P�$���PC(�}�3	/�V�T����^�#Pr�u�s��	 A�'��oCs�G�RN��u��O��h�m�>x	#���B��m��[�̵2�E%Ug�����tH�Ip}������"s�h���D�4d�hݰu�^B^Kad������QAH�c����"���@��8�^g��CV��pzE��.�6�;�Y���Y��0����3$ȼB���h�����N��KmnJ#=�������G(�߷\J��W�Q4V	Y4_o���=R�wx��$���í��l��e��|#_���d�&��SS�/�,9i���r�l���\s��9��߀��j'҂�90Tg~:7J�DW�����B���u��vu�اJ��t� c!���L���`m�e�?�$"=���.�i\ !EH����	��Az�9[��w�����}����I���O���sH�L�z~_@�P�D��\�+@�!Ԁ81�}�`�U̠����\�X��0�6�b�MԲ��y6;f{hEN��.R2��z�����٭s�3/�z�{#��|u�.>}&��@E�_S旈��j).�{� �N2��HB��8U'r���Ո�	������Vy����� A��mUJ�L���'��!&B��/�����mA�Y��G�J��Ė�B�<��^]��@/0|4���j�� ��	t$1��^<�K�4��,���,�,��N����	u�Nos1۴&Z��\�O��;��Ѣ�{Z��R������Y�"E��`�hM�5V���I��S���������]���e��J]�)+��c�'��"�؏Ι���9��Di�J�R��Qw\���%J��e�f��XU�n]��1�(�9�q!��22�x����I��.6N��{#����_92q�Ӥ���7CDa��2^�K�JLr ��ԅ�w�|�r�/8�Xy�D���K�y�k���A�F\�ߐ%��f���X�ڈ}ݕ���w�IlI�0�9�)�u%uU���2��:IT�Ԗ��W�.�`4zy���Cc��3�z-�����XE�lQAʐ���>�s�����`1���U��R�}9�f����g٥;�d�C�
*�ܳ?�J�̣fH�HKX�Yx��]��)��`�Ba[3���N8�.	�4�ģ��WW�+��������ER2
Ʊ�$�t�w��2}�2OR�(_�?�^�Mg���Mk�{ J,������Ct^╕�Zgd�l�D��T�
�Q[�A���7�t0�+B��q��g�Ο�@/|hAM���M�$��{��)��/���+Ƴ��~��!����(�[)ɟ/]��.��M�mh3
,�t���6k6g�(��RM�^���]�����'�c�P�_��a0@��b��ϧz�P�,��'4������g3����m�m�u/Ϥ�I�A�s!ح�`B=٩��j����'��&�nR�LM�V6�Tf�� ���t{�κ�Gu���D���1�6��i,H�ߑgW�C��1T�����g�գ?l��j]R?���������b�"��J:�J�Yˊ��]�b�"��/�;.x�C7�։��
��2ڙO�}��XVC���#D��xex2�7��M<hi�˼xȢ*7������D�?��z���3�w��ݞ��o��AuV�HV�^��}�b�e�K����B�r��]ʰ%7��A����͙xRy��pE��=O�����v�w,S���̾�o�e������ӹR�v�3��!�
��fvޗ�is�lpV�:�� q�WR�t�{ �dNVx����ܪ��Tc��EC��B��.��0s��yX�:���f�Q?iB>��U�|�25�gU8�y�ɾ�Z�K����0��S���T�	v�o�9fӇ�7�VV`^P���S�QLؓ�Υj rd%�'-M�n�KL`\5��= �!�Q-(�����/�-���ԩ�
����r,����E���n�Ԟ�̳��k�j�<��5��'�H�BYsb���&�a�Ѣ���ԓ�s��Fܥ��9�n폔�}�.�P�7&p8&��l�2Mۖ�.kH��-^nbOSJ4��qz�f�>�u7�i���W\P@RDT����hw��:�G1��[�f��Y9Z1�*����"U��ܻo�u��Z+��g�E�f�؀o�r��"������4������|!��]��o*;t{���EZ� dwI��
�*n|e�^!I7x���ߵ.���7�VI�qa���p�O��N�#HP$/�u�,�W�ʵN�}����0�s-хP�#Yؙ��@�u�v;4�) ����>j�s0�2U4��6�!��[�8��k,�)��ϓ�5'�I4���-�^��X�|��8H�ԭG�Ύ;=��J)��Q�㲺�al	)��h���LI�r�ϸ�?��,��vzVU���>���j�����z���v��ʋ�����>�A�#�ԐP{�qoK����&9j���e�|��\&�^Ɯem���"����� �r*t2��_UF�'���u�e���*�[\7��6���?����9t���&W}~��t1�j��L�,gm&)U?�%D��֑au�Y��X�<uL$5H�6G�*3���l�0���b���^�5���jBp��ʞ���x���������e�� \m硾u�󫤷x-��E8����'�����n= ��%=��=P��U,jZO݅;�I��ޱ���H1o��.˧Q-(i4�Z�8ǿ���l�#B=m��;`�2�o��ؚ�~J����}8����3�B��+��Y��;F�]~%��;�o�������Y��S���^V[4H�\��	�j��Ե Ƙ6?��h3jF	�[�4��1譃��l_�5��vqr�h�7���f�v/�Y��9pN���$5�����e��WR�s�ѐ����܏'҃�><�s�����=� -�����a����h.�t�Ѫ������	2Ǯ��s���\v&����@�����.l��Ma�:k_��sqĨ1�v���[,��⒧��d�z<�q�(*þ��H���?��ԇ��Xj�Sͽ����)�b p���H�*&��������b��^o��n[ٟw+q�u�*Nn����<D^�1�G�������w)��|[f��&Xf1�Qb���m�����)������G;�ށ��?�w�Q����G#� �'�+W�&,�b��x�Є>U�82���[g2+�ɪ��d�}j*O< L�c��F�8��`]�Yj�9�{)��g�9�7sN�56����׎�/��c���`��,�I���~�~��)CT5r���%x�\��q;�1
��p�������z�7M���";~��Y]FTFM����|v��Y>�\��
T=�Ͷ�̘F���+���X� (w/��Y�Api��8�=2�@�(��mx���h	
���vŎ�D2Õ���"k�����>Oam3��2�ф?�,�>�� Gw���B���_Wm��>ū���T��uą�Gl�wL��f�]��ve!�:���)T�����4���Ŵ�|��I���u!�>\fCs��1r���9<��[ �������^���V��y�>�����Λ��$A�^M���s<����*��[-��Қ������db���C���ՠ����w��0���X�~0Q2Xb��ǟ��t�<����F�h� ���50*��h!8A@�މ�KvJ�!H���wa�QkN÷�-���4=ow�@_���r���[+-����cӬ�d"���������(��/G4O�p�[>�7c$��賍��j*t���=��u~=#7pG�ן&��aL���*U�o�=~n�I�m�*��WB�wc������z_/X3Gܹ��{[0�$b�E���ol^UW$iThu�GG��wVw�X�j$�D�ɏ2���S���>~O~��!��v�H6X,Yú�DByiV�ܾ��X�9~�Y�c��'�&�^���o��yMD��E�P�D�x���G�X��O���et.�#^�j�Hg�R=�2�d�'�˔�jC��w�v0:kVV ��)2����_D�u��=v�56��Y�
s�+����(X��Y���#���e�1�v9vo.��2r�ڬ�G�lY|�,�
�+��$�e�03V'4����pt��������n@W��!�W3w�u�`���m�D���.��N�Z@5��e����H�~1�Ӛ*/{`qy��ҭ.��~�ޥ+����h����Q���ì��K��Z���VG�1���q,T9�x���"�"�]9��&�x����w��e�(�N�h0���E��g--�ғ)O����?G����N��3/��`q�y�$��ԘIfǻ�H+` _�]�C�⋠us.���Y��t	���&:]���� �-�F?u��S:���G��7F��O>h ���5^�g!jo��"�R>�\�.1}Rh_O��wT(~m��i���o�) �j���\H�������l^Z�AR|[�)�Yn��<�P�z�%A��;�Ķ58q��>@j�}(v��~D�����&�U�&���T�(��'��$l�5�Mע+)�#�j��KG��S���ۯ�(�>��O�48)��ji^ϙ�|/�s��a�c�s�\k�N?�	�O�H)Y���QR"�ąI�iA��V���5{st	����,5��7^cXV�����kb� l��C�'� �H0|.Oh�zx�E�?Xk;���&����|�|EN7���}�xC�,����
���ị	ҔC��Ea�r
������33UѿѠ���h�7���$Y�'R�,S��M����-$��q�2���c$�j	����p,]����v�0��ֆh-m�[7��>45Y�FJw|ӛn������,�*k����)��¯��TΫ���-�\'X�o%����+2��	L�;���ҁ�2^r�e���I:��^�J:���r���(�~����µu��4:Р���&L�9��9?��Lj��?����o��^ٸ��:�Ba�y"� ����.9:~�&�k���#_O��a'(���3G�粓0\;Ei�<�����?��Ж� G�P�T�Hl����#;�H���Ï�,aNL$[���qV���H�t�ml	�G�9���O��b��̰��Q'���7��k	��#]_p�^S�+����7�_�S�CM�����nP�@���a_�A�q��ꅏ�uiV��+�[֡�6��9]mF/zVO>��ef��^i�&���� �6�^e�n�V��;Q�h�Q��`����QL�h��۳(�'�'�䴌��}^k�4X�A-��z2�B1������
� f�{.})i)B\�NO@}�N���W�U�؂q@
�zo۔��V.���nd�%����W��\Hc����
��1�����d���	�(��7�"��j8%%N1�@>v+���%�����D̼̾f͏�Aׁ����qtU�(ڹ0�'a�G���/]�@�e'��C:�&��[!K=Ge����	F�rBP�Ss���ڄ�֖���dm��6@�@�r2��׃Z�Z�c#T�p���lfH�#��Ğl��&"P��ܙ@�MZ6���qw�l^��=S��&��,���řg��]պku���j�s��it�z�&ZP����8?�W�/��RG!��JsB�������n�����hM��]���$�pn䥃�jT��q<�w��G���KM4����??(��Z'�p�ϕ�����?����f���4� YUyo�'���,e�-yf]����RN؄��>(4"�[�ku��BI[�F:�q,Y��]�F �=�d�Re���J��܈HՎ�ЩsrEܠ+�2�)�`�I]|ۓ}3`��-�U��eᳵ^4���/7�0z#z��X٢��B9G3#D����jaz$����1�_�	i��XB�A��$��T���%��������ơ��7��iQA S�i���*�%��+A��`.4�F ���\eWމi�<�2*;Ě6���C$�ND��3����۲�j�W'�Pq�F�}�'CUI� >d�u$�T��l���^��OP_EyuLN��6>�Ay�g��.9�Tgg����Eq��(`�!����x�7����,X����[ؙ���%�"�?���A�SIݢ����"ѸVS�����Xé��&����u���^�����w�ї�-��⣓L�"n�^�mG��|^�I:Cc�{p'4��{���(c"Y"%w��@�0_�g���#�&��9Ԕ�L�7��8Z�ص�JP����U��3������`�J �@W�� V�ޱ_����
(G��Ww�D$����J~l���>?�_)�dX����=�<�q9���ˍlغr�r��f��ݬ�+ƃ�t'߀9��~��ӣ����'l��M"Ƈ����0��TgL�U&O P
�6^U(�,�-~�e<j�$/���Nr�.� ��E�P��ّ�v�zs�n[�!V��E��_��|ʾzC���nH�WRz����]�ٌu��+�s��m �
�	ǂp��;j�wX�t��:�b:��ԟ�y���f�=9E��.�Ѕ��EH��m|��|s�@�6%�{P�0|B�W.�8v�5@�3�_��M���)��l{9�7 lM)�G!���U��A����PڭA���zy�\J�fl�%@�U��
�Z'�s&��`/�T��f��ƴ�G�����%1����<�K]G */L��4�Ɓ�M�-�c	!��$�Y<ן������Yk���C�j����e�	��dN��ۡZC����y��>{��9[�ZN8��?���(�ggh�L5�e���l��j��� �|�&���<�o�2'�J�3+�	�Կ��oꏻ+�wΗ@�s6��Jد^��\�D���Ѥ|1��󽋗��.�;��
�(��{q΄�2{#�~b�IV�6{ �H�����_(�zqM���#�C1ʼ¿��K�L?^��A��ㄢ�}y/�Xf�+�޲K�:�8ju����\�y%/�f�X�}�}j����I9�����˓6R%"}��i~��r��ǆC����$���~�����Ō(c����\�-O9�.��\Q�����݋��ݚI��ڌ�Z� ���}Rmf��� 8��R��zn�0�*����l���f���Ke_Gxjr�����M>&a�d��y�8���
;İ���c�x���L��&?�R_J���j���{���ߓPR�l[_�-�^l��g3�"����z,k���6@	tKm��s�gH^�lX����5��^®Ay4]� t���)I�4?��LM/�*�A���Ө�顒�TVY����Θwĳ��K����)R](����,ϝ�+����m���,�6�I��6k��(��MS;���
�#ڂ���c����U������ƀ�����ZPQݻ���b�'.����3�@�Z���b�ѵ����!E�v`O��v�wj..p�k���*�n�rM�k=6x��a�ꩭ{u�eN{A���E���&ꄂY76� Nv{H��g����l�1�� ж41��~u���]��Ӟ��U��z:��*�"B����k���˗cg]�M"�_a/y�S.	:7�OQ�����R$O����M�+3wDھ3e��7�N^<5� �8R�ȯmW�I�H�D|�T����`�]��w��S����A��>Vh�Ξ|bM��x&�x!��@��R�ҕ[ώ$D��ܞ�΂��p=�����q��$�A�΃��)��D�ۓ���(RK�3��ŷ0<������aՖ�e��gK� >R4����d�������?�����4ə��L���0�t�y�*�:���SQ�Q��.>��`I��?gb�:y�麾�K���ʽ�0S��T�؜�kc�FE���7�x0`K����S�l��`h[�ך�d2��-�6�n�j�`I>��xdo��"Q�*ۺN����-5������2��]fYX�\���C�� ,�`Crk��0)&5.HŸ���YodȘ��J��y��ú��>� ��sk��N�nZ�Wϊ�S���&�K��2����[�)��mn��<SW�ƀ�,`�����bQ$i�ڶ����@�jc=��*�䕿�R֔>��H���d�LZ^᰹��B"�9u��$�"#�Zx�&gߙ�f2�ro����Ji"b���hz46���b��|����XoW�tH�����e q�I̸�
8/|R�b!����O�%օT�7#BqI��Ď]]Śf��#u�n$��T֙��׼d�*~���0�;a��#�OߨM��u^m�4���4�R>��0��\U����G��!�����½k9t~�rx�66)�v��׋&VX�T#�-i����ޜ{��;U2J�7�fgC����.@L)fl�h��]����rª�y{.��G�vFe�U{�>!Xz�+�ͱ�U���i��l��c�5���Ɍ��>��#�I~P(�o��8��#9���
��Ʋ���ќk��e,v�ID����
*��0�,����6��deM{�*�A\7���6+|u?�'��W~h�h��W�*1�_����L�y�m��?:�D��u��\��!���,|�\
Ly�=^��WL���f�,I��c>�^����j�������ؐ�#��(⭸�M0ײԯ I���K���w)x��PE��0�~��o{KLF� �W%��@�j �"�tZ�L�;*A�͊�,�����5���OJ��~�(6g�Z�#��ĔlV��>ٴ6�տSƧ�B��K�<�j�8"�e����B�q��Y2x�F٤I%h���Lo��3��ƦemS�@�ҫ0^[al�\oUPtz���%N s�?=Nph <P	`[*6��xXn����ll g55T!v�7Th���v����Y��,��ʨO589p�A�o݋-��T�~Ɛ����/�'+Z�����s�W��w=<ǳ�%X�>Ua 5à����!�k�A������5>��ˍ���v�s���B���.�FV�:D�:���:�M�u�vGo[9�y���v�7���g�(qD�H���Hg ��3$Ԕ} �jVޠ����5����bM|q�_�*�L��;ڝU.MbV�o�=n��w1*�B�t*�V?�#�"<�:�~����(�wVJO|(�0ɓ]s�6Q���%�w��)k6],*��D����?��QnT�;?5#
M���+�?�,��ފ�>��/�}S7���8�`��R+'���g2}׆E<-6l"�F���8uV�]���f�R)�M&��(�s[���\2�FVv�{E�\�e�2�`qޠ��#�����fJC�����[�?P �>�1w�p�ƅ�l�z�ϵ��C����~��E]KnF����й��-�,�I��
�8&�={Ô�?;F>��+
6�X�
w|�àF�A�����.>�r'ʤ5�m%W������&��T�2����\��)�KdVm�dN2�]?sBE>AecG�3��u�!A_d?]LR˫3p�T��uQ��G�׉L�'���F(؃��!:�[�`o�T��2�c���>��Łq�����#v!iff������r}���f��(�N�a>J��g��H����~��}	���A��ݟ����M~���9eժ���=-��ٚ�P���B?b��C�9��M揚����즕D����{0b��Ǭ�t�~L6'R�34mݍ�b�ʴ���G6@�u�w��JK�����a�$N��k-`W^�i�w���ƿ�b��[ȕډ��c �.d�������d�(V`G���p��vm�cQ�[�ZƵ��Wt���=�}�~��np��k�d�S��a�ʀ���|�"=+���N���Z��u��� �H^/e��f4{��$�pE:�7��`"�vi�%�T���$#����$u�K�\¶ԕ���~�X��.͇�#�6��Bç&ZB��	���%5,~�P�c͠�Ӕ���	�\��y����BZ�P��'����*'�����@�R����>�j,;��u2T?q����x��j��w�9�v�Mp�%P �5]2^/��{D�I�[�"��V�IE������d�<e�BYB�hp������1!��2�l��G5�G';)Y)|�WY�+������33�x�4���k���@?����F�@D@hᮥx3�Ҹ�-�˅@0D����UNb@"/em�u51�5M���{m>6����F�߰L�2����Ëh��/N��%q-�A��K�O��Z��^���>L�9x�x���� q��w�����h��\Ge�ŨNC��������;z�����OK,�lۋ��NO�/3<`#`�UP&}���I�F�u�� ,�������	�u n>���a��͙Q:/���|�"K�U㍁uc*�:��G�t�FG�Ok�fз]Aˋ�g.b�Wδ��m�\�G(}ߞ9O��T�����0g��$�)����T��\�Mz�ҏ�9����6�hiB)��n���~z��ƿ�i���9h���g��P'��B�c�E��k�W�����UGE���<��;�t��56x��X���$�jn�K��� k)�(O�oR���t��|4�8� �jֶ�Ϧ�l|�����c�PZ��K�ᡸ�;�	��2H67�:D�Ro(��r��iθ�V��J5H�����io����O�cEW��W�k���l_ԍf�s-!�0)m�O��4x��̳�kh�n�x�;��s|��YE��j�F��x0瞧B2
��i���-�*�E��
��w���=�F����E�Qo!7��G�Ѯ�t],@2�M(�@K3�$��eqRV����� ���@,J�ђ8j�Hqw��nۆ�m�h�����>�:���J���Ȍ��ł=��Rk�<�ւ���H�A5�`��Ӊ"$X�Р%��8������j��Tr�=�����:2,�Ϻ��8@r�?��~$@Ƈ�jd�%�:=Uj��Y�L7��8l��oɵt���$F#��g��%��G�=ae��"��Y��L�9�;F&
�����M=O�\�a�e�c}�34P� +�;r��<��;�<K���� �1��DEHY��d.M;r��卙�ML1�t���V;�H��m���tF9v�x�E�o� y<ڞ���k���@�P@.pQ������xش��S	+��n��1]��mzk�.%�Ai�����1�"xF�^��H|�kb��;��mr/V���)�w�y���*���G�C���ߖ��-{VPa;^�h�t�?m��G�Q٠\�3(��������w'}��]��.r��B^�C��<5
\����}��B�ÖO-_5N=WW"g�O�%
d)o��R6 ���|d���]M�W'p�\�ĩ;%�sB1P�f�8�Ndp�V	�L'�����2-�W��2��1��+vx����V�������j���4��N,��~��@��~���9���R] �}r9����	&�C>�=�\d���	��r��S��!壋}�#]'��'ٶ��s�c�@��r�Wfא�)��$#^�6�]����0�P�:�k�@�P�ʙ��Z��o���q��^� �= �&c}����=��ު�Lkb����s�(t�H&�ev�{;8�qW��	�?K!�so���`f���v=MFt�Y�]p�Xj��{q	ea�r,d���M�`~i,f_ �')ب����J3�?����,U�0Ϫ4}��U�>'�?,2zy��P�����p,�=��4L�����opI��R���m0
umFMs�QiR�A��w���U�z�*� sv��l@�c���M��L���^�`ߓ`-'69�r�յ�e�d�*�����wz��2�o�B�Du#Q6&��wzh��ӹކ��+�6{���Bf\��1FT�2��r_;�t}��R4���h�%�ֈ� xiix�n*h-K��Q�A]�^.a� ����U	W�k<io`��_˙;�]��>�:CQnD\=9��_�ۿ�{�'^�3P^$��
�C�%Z��2���CT��/A}^G�ZPLB�u���c*:AFK��I�t�a��T�2�����-��[�ǰ�x�&Ϫ�r�*.Ƽ�R[%'2F%o��lU��`IJ����e��eK���n,Y�1w��# u{p�^%����Ǜ�D5@�:?����"�A�������5^Ai Cp�%p�⩏�\�q�Y��J��}�0,�\�ݴ�3Sƅ��fƙ9K�����e��J}�����<]�����9ɁJmM�Wr!�V#$�_��7��:��w�Qa$=�Q�G��l{�k����_Vrnd%5�-���I��9�[�D�l�<�v2������yn���c�'�>I9���~�a'��ي'�T�[�����O������Da���� =���×�U���N�e�T�$<�����!.\�_ �
|Eb����tC�z��[�b�6hв�տiuU��y�:��Hv"wzX��jP\�"��+�ܲ�Z����ƀǯ�̫�_�X
�O���"b�Z|Ԍ"3y*яf�PE��.,/я�q��?�6�4so��Ï�{}��|�t.�;!��@�>�_�栈��)H�{fby 9�ʹ�%���RU�������zW'�Σ
 D%yi�C��ˌ�2�.U��.2��'�^�&\}/������3��G����wG��
�<��g]�~a/yм4�<O�D���:�	�a�q��<�}}�N�%Ά#���hؖק����8	el�N	V
ێ=Z����d���Cܖ�5�{!H���r>ǧ����W�   �   rec�jS>F�Z}�I�CAzmi ��H��%R7W�L��$?��h�z�piS��?)��K(��9�Հ�.!Q����ن
�4��[*�M���i��!{��⟀���4�M;0�&�?�!����P#GD�PU�d��((����g�H�4fl����BL�""�'93�[�pFD��/D�;0��6nJtk!�"?v΃#L(�� �<��Hڴo
Dp�F�<�h���DI�2��=-@b���EE�;C8��S�V_?a�'N�(GH��Q}�O?�i��Q)Hߢ�	�O�&lbT��%�� '��rw�W�%�r�OH�r.����ٰ^�`�0V��?�,�QF����>6^�u�ѵi�Zi@�`f>5�!�!hR���<) B�,V::�Xp��_�x�C�#U"?�r*u0�De��5¥�|��O;/��A*��	vYR�KO�-��s�"���.�!���D�$��~�Co�����>��;��E#&*L�#AhMJ�8M�I�}H�#rc'��/r60ˢ��'|Q�Se���
@е�]�i��%(C�@}�0O�������1O�rp�
&�M���'�0��&��^O�q!��T�\6#<��a4?A��NtI<�G�z��5C�LyO�S�'��u�?��KŨN��PAti�;��ase/S�4��#<1��(�3,��F)9F�l�A`�Y<�DIUM�l�1OrE���dX.��H��AӇ��MH�ܠPK�4w�����se*#<)pN3��,g���Z�Xd4��hA�(#L��g��+�V<�7��=��P���S���!Jn��N����*�
�� Uc����B/B�� 0��� )�2H�<���*
���'�Ș4d����O���1
@
q�*�A�BdP��=Q�p��7�|r9�b��y��H�.��(p�!!7�ڝ�^�u}B���"OzpYB�  �@�?9��'��@ ��                                                                                                                                                                                                                                                                                                      