MPQ    x    h�  h                                                                                 �gI=��	�#�V�)Qv�@>A?<#�Q��� oс֬9�`��v\h�2�`aՀX�G��u�г�,�6k�M3ɗɥ���
�m����A�bꆜ�S�$M�z�k�ws����s0�z������a��@Yޠ�{ch�N�}�
!X�9	e�ɱ*��D�q���+A#����oǸ�c[E���y�:̿�vp��%Fs3C��+{���ݺ;+���g��^V[�B9Fy1�_�Sn	�& @��Ag�EXɯ�~g;�yIbi2ܒ�TX��G=���$��)��q(N��-�G�_��S��a�����?<�3��X�	��+�nc��G��j\f���?�~?�0�!7����0v��B�} .s��G����4�&���͍(�!��+�|�d}���2񜮱I������%� �/��,)���E����_�w�@��ˌz��$G���U�г�X;ho,R�¡�������S��~Y+��eE'�x�t%W��D����J�MO�۾������j�X2�(|b7լ;� ����p�d����c�fϦP'-���7GS����M��3%��uԡ��f�X@b=.�#P��wL��k��aə%L�}*���%���B�q�������V�匐<�2w��T��k���%}���z�r��)�xl[]U�{�:����9��(�1�$+���V��q�i����P^��6^I���犪���U��ڲ���qOj��S̗Ut����j�J�����E�5=\S}�f��Ct�iv ����W"k�WRIg�&A��@cW��6+@��h�!T��qiwN%�Y�z%�ީh��WX�\��v~-8����b�"�ʸ^I�-u�+h�Oc��;Z��v�P�BC2`}!�=�O;�!��]x�:{�ǃǗ`�AO�1�|L�I!�@�m�/N*?���o��>����k6w�$�[V�;`{�!���< p��*g��1��r��%���n�y�h��COVoW�'� 	�P���vnBx4L��ef^C�ׄ��˓�$F��-"�$�L�U�t��Ku2	6�h8̄�hJ�-�|х���俧�7h�xzў��ǁ�GVft�Ê;���&t�w���s�Qu�='ˢ���6W�k��V��H?��,1�XV��PMK5�`��\E��˷ϳ�Jr��D�Òi\�Ҥ�RBb��S��]ɻץNo���LY�ȟI0�_���x���/Ct���s����m<;�cN��yt�%l�H8إ34����Iu�A�y�����n�*���Y�{)�k�⯏�q�?�$چ�Z@Y�uTf����e��F�|�Z�}�:�ET��cv^n��t��6���{�ѥY��QQ[s` ?FV5�<�1�s�ς�����?il����k x%g�w�ř�=w"a��2ɷn��t�;���s]v������g��䁿�S��s1�tt)�g=K�d$ɹ���	'2��"�_{�A���԰�P�A?��?�z*�s�9����
n��FLٌ���*8K��w������*^�P�+/XT	�	i��#Ng���YӲU�5��O����7}������H(�|���uce��vk0�����P}���1���#aL�?���+�'ۄ�H�8ٛ}t���}����չ�dnW������"�o�h�C �S���MT^�ł��g�~��)Z��}�����'���b�]�l-p{�l��ۚ"���!��+��[�����|b�M�B�/.��瘛�o��\Ps�x^��Z6=%M�m���]?$o���\�"}C_Z�L�/ӄ�h5�2�H��D�~�\}6��ԏ�ÿī�c�~��w:8cli��m�!��&��Ĩ4@���c5џ����M�u�����j�Y���U��Vs���"�O2o� [^H�LK�&�i��aacMԃ���V�_��v�A�\8߳�͗�R�y!Y�8���Vp�w�V��Mֱ��Y��B�=~�_�-�XK���tN咹����B�Ҳ�c��A���9��[,[�.���� 3�=|���o��{Q�cl�7��`Q��OD�z�g�W%��� t*�VA��3>|#-��[v~�����Z����`9;҃J��$�9�3����m�b����YiLG0�)�_�?gL8Tr�'��Å�%��5/ş���� R.5�ݒޔ��\�3,G@�l�¨�����G��*����r�#��޲ܻ�+�.�ed�g��<j�
h�ՔO�g_iV��]�
��q��wfrR��u��%������l�>m�܎�z�?|��&띚������22��D$�ȵ�r��\�Q��?����--��Llgt��q$�u�"5�����O%�O��ާRT�j�ëUi���jEfOBXEaT�
�Ïs��!����,��'����JՃ�yE9�����f��i�7D�'��;g��3�4�X�'��zX�l����e�y���$�}����I0��W,�H���FyVR�q��ӓ�{�f�0"�HQA�-��g�Gє�����m���Fׇi%��3~�]U�}���R��ix0=b�$[C@�S({��Yf�jDǸs���Q�uI��@k�a�>:�����V)E�ǃZ���a�D���޴p��G_�(�t��5�S�בu�*�0:fVjw�I3�&k1Y��+o��)�r�SK�T�)ؒ�!�GC��/p\ҏ$QȊ�
~mW�W9(e��&H��7}÷���9��p�+n�x>Kf��y8�Q��C����Eθ�l����#�aE%B{�i�c�S�Λ����d��w��l/m&:͟��V�� H"�m��k�W�e�/{�HR��w���ڮ}b����Q��1|��w��y`�Y��M���,��o���iHO0E��D�y��|�$+��ۆ�UGEg�����l_Fh���y(�L�.��n�~�f��YUE�he�Ad/ w��.@�ֶϩQ� �@��A2mZ��
��XC'�8�X�u�.àT�1��ՒK�V���l��p_37=���)�Y��uYZ��!Q4����-�Y�@9��<~Fw�E�;�r�Q��;��v�S_2��@a�&C�u�1�ڔ����M,Fbި(Ρ����0�]m�'Q<��b�"��n��M	��k̽����L��`7I�<g�>�3a��9YYb�{>Y�N��L
���9lW�$�Ώd��q�n��M7��%o��͡a�E����B�%:���v��"%��]CΠ{���U���X��3�y[x
�9]1i8SI��&[m���;�@�ׯ�sYg�H�I}����X�0�GxV�ѤNy�Q�qO�N�`����:�S"ܲ�&���^Ě�(3�5-��]	�K+\a%�ȕ��rp郻c���d?�$:!Rb��}��0Q�>��}����۪�h��b�T&�B��H���;�+@���h�ؑn�	�7�����w#��>��6&�����_a[�2!q�.���a����E�U$���S0�o��A�\�S��­����Jf;�e�Sx���t���U����`�Ȕ�ۙٗ��hjo�a�#�70�������^�du)��>{.����-�ʥ��FG���^�N������Y�ۓ�6=�d�P�L�绯���@̑�P����B�dB�h�q��#|Ǎ�:� ;<����Fx��'fN˴}����rh5k���]���{u�0�ɮ{�3k(䳦$�St���q��i0����^����&�I�X���G͐��!$�i}�L�!��>��P�Uo���qJz�v���G5�� SX羋,��X �w���;k{�I�@�Ap�c2�+6f3u�I�!O5P�̊�w	>,Y�-�$�h�y�W��ŵ�<-3))�R��"�n�^5d!��2+CcM��ųk0��ԫpgC�:!/�w;u�rTʢ��������O�Ǣ1�mu��5�@z�/�I��H&��H��r����6���Ey6�+;��ڝ���7���Jojga���9���t�|��m���>��o�R�'��	��ll��ɮe��ҿ��e��+4�ʰ��2��02��?uͻ��c> ��-�����Ѡ=��_K�c�W��zl���RG�VZ�~���JtN_��4@ߌ�+=�S0��%uW?���x��c����Rس3Sl�N1M�(�`�NG\�D(�r��e�[����me7��R���N�p�:�`�8�5�L�r��z�J�����؍�,/�(�K-�����m�=@�>��ô@%�8�m�4WK0���2K�y'ě��n˞w*V�bY���Ɩ��Jɓ�Z��$�r/�5������[��e~-�JZ��r�Ux�EϋzcQ�U�"5F�/��4,ک{�%�Y��Q��s;�F��E���1~g<��S�<��i�k�[��x���g�;P�4a�=r�G�s��2�2Jnڰ���b;lGs�Ee�`���b9Q�܈oS@�E1� �)w_K��_���_2I	"�T��o_6P�A���+ceP��?�l��n���
)��Fg;0���<K����Y��j���+��	�Vn��s#)g^�4U ����+#k78)�����p(�'x"#bu�20�q�p�i&������F��l#�]܅ڼ�a�������O���݆��7��A"��{OWR��B��=�J���} q�0�W�5M�l~�}d�g�̺�5����~����}��)��]#�Kpv��laEK�U�����A��_��6 ���Ub*2�=��/�3S�S��Ɋt�\�q�S�Ǖ~�%��I����?��NJ�=�s}��ϛ'KNӿ	R5t�H�DHdk�����d�>S̫�f�~�H�:ӈ�i�(��ǿm*���#4��u�>�!��SC��z7u�1aj�~���y�U��sjlի]S��j� V��7�T��
�i��a��4�d�FV�����A͖d������y<�7�E��1�w)���~3MѶ��<B:ܪ~���-Vc�K�y��
��-�����a�-��c�ЦA��
9�C�[`�.�i��<�>����]�!o���Q�`��}�`,W�OE��r%��[&���7V\u.�)�#�[����'�U#��,��;��o�|�6p�3�"G�� ����|	鏴�G��J)����8/#�'ݑ5�yq�0�ڟ
h��Er�.!ޚ����b��3gl��i��q�3��oϕ��h����@e����|�ƿ�`�hg�
%��e��v:1�B�9]<���l��w�����ڀ�X��u����%��m�܉�uu�|BG��X8�����*7�,���0r��>�L�?zM �fVD���Hl�7�L�%װ��5e���qXO�S�q̿��}���>��0�����E��X�TY�u�J��<�v�u腻⢼�!&Jp/�y@&��7ϰ0e���DL��g���&���5��A�'G-ez�߶���e]���X.���3�I&0���,xL�Dմyq)�qE�8����fGD�"Q�mQ<�_��<X�h�*sۘ��@��uE���}]P�r��IR��V��%#=��l[f�������a����sF96Q��I�k�l�>uc�9׺)@����Z�\�a�Ǟ�Y�Lp���_*T�$`5������*o��fq�e�13���kl�dͳ.y�t����KPvp)��!��`C[����%�*|�L
�e�8W�E�9C�ȗ��H�O�7�U!�X��ǯ�j$)͆>f�W��J/,U�CRT'�T�����Ѵ�#b$�@\/��=U>�v��v �#w&�_d�w���/(t��F��J� #��N��m�*S�{�򇲴���S�c��Ō�x�f@��}�K����E�C���{��ٔ���"��()��.WĂ$`F�{m�O��n�3��RB|�a�e����)FE����q_�%����g�2�,Ci�YT�59�U�Ah`�7d��ӝ3��R��
��t�|�Z-�%����'*����IJ�Ti��аLʿ���c	��k��7�(Ǌ�D��t��u�������3�!-ga�@4�V<٠ ����V	܁̍���v�^62>\�a��	��1ѷ��1�$�,��=���?� �˥�m����b`�e���M��k�#��9�(���0��&LañZY�C�{j�N0�O
W�=9�����2���q�wS!z��^�}o��<��E{�5睼k:BY�v���%<B�CZ5{G:��.h��C���[3� 98��1��S$�&����w0�;H��6�Tg��.I��܈�PX��ZG�����0�����n�,M.N����׶�S]?Ƶ���߷�����3u�e�8�	���+7tW����r�~������?K8a!m����0,F�y�}6O����^��0��R�&��f���"�פ+{�W��tĠ�(�dN!�#0�9G����R7l�y*Ȓќ���?=_��n�Յ�I?��p1�����F�)U�s��NEo⚚� ��,&���Cˢ2L��e{�"xϸKt�������Ƨ�C�-�t�f���j
�I��c7��c�,�.k�d����;F���-P6ѥ�Y2G	E����i�I�k�m�uĬ�ά=d��P�G�LZe�j�[� �s�y��1&�}n�BKa�qz��b��H�é	�<x5���L����.|}�e<8�Br#�p���~]K�;{P�8���U>(�U�$�45����q��ei��W�Ҙ�^���`�I�{��@�1�e���&�ѐ'���y݉�4Uj �n�GJ5����53b�S3TG�B4l�Mhl �z��o��k6�I���A��c��6�FA��=a!Jn�'�w�v�Y��e�h�<�W�ܢ�2"�-.��ϭ�"O2^P��#��+�vc���N��O��T,C�ݛ!J>�3a;P3�?���=�p���g���O��X1��?j�@U��/Ĉύ�LJ�BΧ�M�p�6�������;�W�A�2jI���m"Q�� A񂚟����rt�����9Oo�P'`}�	��� ���)�e�����C �Қ1�������,=�uh�	�^d�L�{ѻ�u���l��}���D
z�I��CnGg��9��3�ut�D������W!=]�յ���W��E����~.�"�ֳ�2뉟�M�<�`��/\��!�-<��$H�:��H��H�Rx?��I7��R���PW5LOJ��U�U�ժ�&����//�̠�u���8um2`�����%�8�8�U�4�2᣿��Muy�xQ��8�nW*�Z�Y����!�j�'��u��$+��� �����ey��`�\ZH�̖px]EJ��c,$��]����}qB�{Y�rY"pOQ�ws<�F��'r�1y{��8�����?i�A���~�x�|4g	 ����V=m�j��y<2���n�q�j��;G�cs�4��z��]�t�7rS���1���)���K�#��u��s 	��W+_���AיԦ�|P��?/r띰c�i3��ELJ
��hF��{��v�j�pKQ�ɭ4�~�� 2�Zm+���	��;
��#�;�op��������_~ �7�i�T&�~��(q�x]I|u� ��l�������=�����^^��#׎j�u6��͔ݑ~W�5��Lzّ@����?�M��$��|�lW�����\�Xn�^ L�~�==M��n�xf|gKႺ�����-��	����R�d��]��pq�l�������q�!2��"h�3mAb�6f�8/������ɥN�\F,�.�w���W%�lޝ�V�?��*�	XZ�X|�}9�ü��|�5��H���D�Q��Ҏ���#������:~!�`:n�pi��o#��(N���)46�6����=��+�u��"qV�j{-;� �U�	}sE姫���h�5 Q\��	��D�iǃ�aYV�?ͅV~d�A����i��J��yW�.%ʈ�wd��ՌpIM�۱�gB�+~�͘-э�K���>����R��̴�q�cn��A��9��[�`.*F�׏��9����otc�Q�},�->�`'�O�����e%��ZǶk(w�
Vw}_)54#�D[��1�|�Pt�̇!0;H[�o����3�H)c'�
�w%M��{G��%))�Z�5��8
�w'~[���T�+�,�e.B� ].<��݈�n�=4�3�l��uh��2L����*����h�@���(�1�a	a�[>ggn���)�۔E���}�~]�S��g(�w��ʒ�	㨵�L�Ӡ�}`�jm�<�p��|�������*d>�(CE��Sg�>�&r2���Gv?���!���/-l]��'������5 ����O��,������`풫Ez�%@�E��X�T��
�J�W��������\LJ�y;eD�K�k���D}�1�B�Z�a4�1l(��Kp'�v�z�S7���e��~�'�� ]%�z0�X�,ӑO���&y� �q��)����f��?"��+Q7��ﺵ.���?�,J���Иe�ڇ���iM�]KT$�p�(Rx�����=XO�[��4������\����s�Q���I���k[��>��N��$);���9{�<-a�jN����p�i_e����5�ˇ�G��**~-f�f��@F3|�k�q��NR�����(jFK��)e�!x` C6����
�Gl�����Wy�9^���EH�&�7����JZ�&7�$�>���o}6׏C�ť�����Ӵ_�E#�[���_�8���#?٪�F��Z'�wO�4/���\�L� ��$���mDe��vg���ڥL�~���e��{v:}����-6����6_8ٯ���O���W�i@���p�v��O�k�UB��8�|�W��@mF�&�E����껲_�䃲o���^~��7/�4؟�p8�UI��h[D�d���XX����GJ��>@��&Z� ���B�'�A����V�d�T�&�Ћ&Y�� c��L�f�7�w��AƏ�@uO�6��:��n�~-��@/�|<4
���2�q��G����"�v�a2��a�Ҭ�+�зP&�!�b,<���c��z���f�m�i��R�b���� �M�=hk����t3i�M	����a��YOE\{��^Nk
�r�9�ّ���V�ڹiq���C�9��o0m�׾�Ev�����:�ըv���%���C5�[{��݋�:���j��s�[���9S�1_��S�>�&�'��E{6�ȯ��pglN�I��"��PX��`G�&_�P��
��A��jN����vP^�
�S��-�\�_���,�P��30g���	wl2+���>��;�l�y��P�?l!���s�[0$����}����c.��t���&O�>:b�-3+�=Ӎ5���ί����zm	�T���,-kִ�U�l3�ũ�_����~�d�͌� XzaS����UZu��Iz*o=o���_6�G}��/�}�]ܥOe�xʸTt6���ˤ&��鄹�\�O#f�2��j��}�7��W�Q���I�ydk������W�V-�x�����Gd�����ք��Ƶ�PO��	�<=��HPΨ1L��]�%���v�}���v�zgІ�_�B�y�qu���YK���6��<��[�w�ϧ5 ���{}�\,��1r�X:�ɗ|]ƙ�{+~�?�{��h(�\$<6֓��q�Li&?���x^F�g/�XI�U������+`��n��b����$�gUeX���>J�2Ն�r5�?�S���}\6��{ ����~.k�`�I�*�Af�8c���6�ya�؇!E�g����w�"Y(k��٘h��W	���'-){`���"
�^k���P+�bc�h���,%�	ӟ�aW�CcL�!e�T�j;+l�z�(��l?���q��OI��1-��ĺ�j@0��/��Ս~��\�O���+�86�C�d��;Z-��GR�-Op� Xq�`��(7���VvР�菢9��4��oh��'�	:�=�b����9��We7���ȕ�����UW�-e&�����1dg�$u�7�Y������^6��֭A�U±�ȸc��گz�W���T�Gg����ݳ�NH�t[��}�����=�ē���FW�����p晹���� ��T���KMpQ`�|T\V1���d&���|���L�#�]��j�R�.�D��n}n�քx�k�L�A1�0�P�mI�� ��lR/T����#���m��N�����*|{%=�d8�]�4:��z�ށh�8y���uenA/�*�:Yؔ��|ێ�������$���|�&���et:��4�ZՊ����EŲTc�t���E�e�}��ʠ{-�Y={Q�<s�y�F��M1t��ϓI����5i�7j�Q8�x�eDgD$��jX=h���)X{2Mf�nS��;"&PsD�Ֆq��X���{�S���1y�)��Kdb`շAڕ�o	�O��_�_��qA�P!�!x Py�&?j�ߝK0\d����(
�(F�_o�\@E��K����(\��K��a�v+`y8	�P���5#��h���V�&D#���pٵ7���/���Z(L����
u4.��gN��)���72V%�<%��ox�#������Yɔ8��MD��W�R��a?�Έ4����c�w	�W���g�sAل�x� '���ͤM%��s��g�B�Z�����t� â����Y�]Y9�plm�l>���	����)��$���c`�n�Ab`[v�3�&/?����#��H3\�iq�	ŕ�o3%�*����?5�ْą��sa�}����Z{�5!5�¼H� *D�^e��G����H�4ڟ��~\e�:	4�i���~(���S�z?4�����s�Q�����u�� ̹�j6�!� �XU�rRs ~*�ӛ��� L�헧�W�i��a�
ڃ�VR=�
�A�j���n����yrm^�$���w����'��M� �j�B���~�4�-L�'Kk���y�x�c����s���c)�8A��9|N�[���.P
��rw~�n2��	o/�Q׺8�%`��O����8&1%�F���2�AV��x�`r#� H['���̂��K�����;�F��,=�3h��Vd��3&�ra͏j;Ga�)D����Ks8���'S�5�Q�p�&亟��򻵈.W����M�Ћ3�,@�=t���������(� ���n��&�c�ښ�r.�V��g�������)��C7������]r(Z�b��wwH��M`$�f�k:�{3N��Nm�;��k��|�K���a�E�%��{�՛��yqr�1��Bt�?0�o����5��l؞����&Fh5������O6��瓗��3��ۻ�����`��E7q�X��T�?���!�r3ݙk���������J��{y6�����&$Y��T�D����������¦��u�'��az��r���eS���Yv�.�z��G0�M,.&S����y�7�q;���c��f�.�"�)�Q2c��u§xqK�GL3 �q�@Ť�v"���]Fߑ��sGR3�
���`=��a[ԅ'��R�P�WY�U��s��aQ�I�,k6�<>�1��o�k)6��ǔ��҇a�-�O�pk_�_�Ug�E��5���עW�*�Tf��[��3W��k�-���5�
\�܃ `K�E))�q!��Cg�!R��`�LB�ȟbpW4��9y�̇��H��7.�Е��u�i��#���>�S������x�C��v��sθ��q��ɦ#�	ev����X��M�^'ƪY6��U
�w� �/�oS;���q ٗ�ě�m߿=�q0�ho��`e�4�ł�>�t���t.}3�v���"���n��'��������ޤƤI��Z���qթOA/nqn��>�|!S�f��a2`E8*���/_WӢ�*G��O�"LA�|��W�U��hV7d@��8�'�թ©��э���PcZc�ĉ��;'��B߉�����T_�&�f ��6�����aO 7N烊���ƪ<�u��t��ߙ˩/-�Џ@*�^<��3�=p���#���%��r]vH��2t��a��+���0��~�<�,�����^̗�>=��nm�:�MC"bֵ?���-Mz�k]O񣯔U^ց���.��oia�MY�f�{��N�nr
�f�9�@��5;����q�)3<���ok���rEq%��S�:�r}v��"%2�eCc�{��&������D�[�!K9n91ک�Sڐ�&���y�1����i�g'tI��m�~�XwǖG)�T��Ov�z�b3I��DN������˲�S�e��ˏ��S^ī�3�/���	�O�+���y@`��r_�t�2��P?��;!�c-���0�!��f�}l���W�y����&.�չ����+����ܠ�nO�k45צ�oi�����嘆����3_rWVc�[�7I�f0EU`���sU���Dϸo�cL߭�b�`���d�Xf��e���x���t�,ㆯ���K��9%7�*x��m�j@wA�hU7A��8I�d��d����fϒ}-��g��G�̚�#֟E|�a�+���D�m=�m�P�)�L�Y��Po���i���U�
��p7B��qp�%#Ǿ!©Q�<n�U�R��pfV�}�sX��r�Ȯ��]A��{*��z�9���(��@$�WW�BS'q.g�i��B��&^� �3bIԵ���Οx�ˁF/�� ��c�V�+ݿ�2U`���$�TJ����1n5)=wS�苸�4��B ��t�%!k�N�I�ϤA�#yc�K6�����!@�=�ݒ�w:H�YC���lkhp"�WDy��hMr-$T��c�:"�`^�uZ/�+Խ�c���ń�C�w�Լz�C�J!��/)�g;���n!�shF�����!�O�1H��53�@�S/:g���F�`�� ���>f6�>%�$��Q�;L�ĝ�۰(T�[�t����4O��x��Q*E�Z}���K��/�To�`x'�Ҿ	U���C�˛8J�e�<���0������Hb��������su��=�Tń>^�����Э������z=�򩳅2G����9��i�t��]�X��=��=��i����WP���B̲�w�wW�����M���`�C�\��Tˣ�ԩ�V��0�^�����A�R����?;��Njב�_8LEY��;�KO�\�ȍ��/����|d��)@m((��U��ei7%�A�8ą;4ha��5��)y��p�a� n|'�*':�YӇX��-�{B���=u$��Ɵ(�a�!�,y�eo���Z������CE@��c�i����s� �mo�'s�{��OYX��Q��s���FBڧ�E�1o���R�m�i�ML���x�ngHw��=c�d߄Vz20�n+T�`�;��sIs��1���S�����SqK15e')�eNK?����0W7	F��y_g��A(�Ԝ2PPT�M?����m_K��*'
Z��F�!��aT >jK�[�j����������+o�	�. I#�&������x��]4��7iKpJd�t�4('����u�[5�b/�z��⳿(M�7ͷ�J.�#MQC��&'�ᔓ������	]ه�8�<���ð�Z�X�r�[Wc:Us�6񎚌�T�� Ê�,�M�XW�n�|gď�M]�����x��}B�����]�xpgzOlr�5ۆAع�j�7����h���Vb���.��/�YV��[��bR\<�s�����FC%��/��|_?��ȒӴΎfF}/A�����p�5E�XHӎIDY�r�H ����V���k�Z/_~�#:��Ui���ـ����D�0U]4,ݰϬt��O����bu���'=�j�ꬦ;lAUw�Ss�6]�p>�� G�HF��i��kaO���ttV��U��A��Hܗ���y�	$D����#w�l��³�M����Bk+~�g-�BDKFGV���Y��k���f�>�<c���A
�99��[�.�.�
z���i�nG^o�aQ��#�`�& O0
�Ә�%���lV]�,�V��y��#�ۻ[b�q�g` �Fv�=b';��������3C����1��ZY�m�i��+GI�)_K�+-�8���'��Å�3��!����v�x.r���~�x��3d�ؒn����D����/�;��^� �]�ޞ%x���s�Q��g$NuVlYԢ �;���!��E]q�]�w��+��z?W̵�G<�V�N�TgmQ�ˀf|S�����`����������rh���=��?��������PO�lSBM�ݯ��a�g56�筡�O����������V�����q��E�\XU�Tj�{.����̙�4��s}���4JA�y1C��T���My�յDsy���ʎ��2Mg9}��^'Xi�zD����h�eΏo�45�i5�[��0�b�,��V�u4y�n�q����>cf�Ӟ""vpQ-Cd�pTv�3<{�bn\�C��ڞ�U&_埜�]A���&~�R�KK���=N�[�Ej�?U���R��܌sw{Q��FI��SkMC>&���
 �)1*���P��a����8]pFu�_�&O�୽5�í����*�K�f����C�32j�k
�̈́���3��޶9K��U)D��!n�#C��\9����
=�@�vC�W��9�5���Hy4�7i��)z���/Z4�>���eB��:�C�<�%T��%��(#�,�j<�Uό �/��E��P2wc�/Y�9t�B� ��|���mz:w�l㘇��.�����N��#�OO�}Μ␅?�TSj��ƙ��G\�E�����r���l9�O��˿���d�|�
��~��f{E��q����_�ၲ� ��`����?��{UhhQAd�E[����B�R�=)�ˬ���-��Z�#H���1';���D�H����Tڛ�A:��B�s4�n�\�|7�v���T���xuE�^�������-88@%H�<�o���u0���ȁ=O���v�@�2t3a�������;�W�,2P䨔ye�������m�+4�S3b��r��&�M�
.k8y����~g7Aj�*�ma̮YE��{�\�N���
(z�9�ǼאqߏP�qS������ԏo�{o���Elw6�:s/6v�@�%�h@C�)�{������H��/��[di�9�A=1U�S��&Gb��H��,�*�GQg��LI��`���UXR��Gdw~��� Z�E�]�N�m�l��z�S)��������k�/�3�h��	mS�+�l���1�qJ�op���?|3�!�NO�i/0�?�*@}���k"�Ԋ��N��&I���4Me�h��+,��kW=��M��u)^�`�*��՝�2��*�풢�����t_�@�����,��_�0a��mvU����?D�o�w��H)�}�P�G�30�R�eLF�x�;t�S��A�$��I���������gjێQ�sh7�� ���J�R"da�A�:n�͘-!^���{G�F�JQ�ֺ���]
�����=5[�P��DLkFջ�c��[P��*��03Ն.�PB\qkw�s��yx7�l3�<�{�-
觫X��#}���I�OrT����P]��J{��2���&.�(���$򘸓���qIkRi.ڋc��^�R�e��IςB�Q��3��a_y�����E��Z��U[h���JfĆLH>5�Z�S�Z��g�W� �C����!kg\CI�8A\��c�ð6R@��m]!;-�8�w��Y^�_� *hKEeW����-M�Ͼ�"�=T^���-+���c9[U�nz��:���;Cى�!�p3���;�=���������'�O��1cr�İ�@��/u_������3��+��x6��o�H� �;��P�(ܰ#y2���xS�u�O����h,���2�o�`�*�ZoP<'�� 	p��X�f��-s
�em|ݾ�6T���%c���t1ۜ���>Zu9��O�i�]����������K���~�p�CgWz�r;��֎GX��j���)t��3�x�z=.�W��ՈW�4��Ҙ��U���ڳ�֦�:�MR7�`�*R\���^hG�����s��ٔĖ�8,RI{��:��$@F�L�H���L��m�����Q��-	�~Fi/
��7Y�D�qm�����'�àv%s�o8��C4è����.����y��<O�n�?+*�Y�YΚ��2���6 ƑƲ�$�ˠ��$��Ģ���ej�_qO�ZyF3��8�E�Y�c�<T�.���U��;�{���Ys�Q�y}s�U�F}FC��1jw��I��(si�V�G�xd�tg���Š�=^<��t92�=nFu��&�;ح�s��	�̾��N��H�S,�v1Pq�)�� K@�KL����v	;�h((_"�gA(��P/ӄ?�A��)Z��V�E
�F�O���/K�K��>���YJ+քz	5�T{�(#���� ���\��'���7$�^e���N(|�uj�|�]0L���K�n�h|R�2��%�#�⍅F�Ø�������M�!�����!���L����m-W��Y."����ϑ_ ��H�C�KM[�O�i,�g\e����w��j`��X���]�wpb�-lͶ��A���m2��i�ӢG���Db�_�)�$/�PB�?�����\�D"ؿ�aǁ߆%T{�}?�?����:A�Ω��}�	�����ӫ�@5��H�ED��߳���L�*�#�5�~�%:?_�i�O-4�`�Yy��KP�4�b°����8��T��u���j��ۦVRRU�s�@�Id|9�� Bɪ���ͱBi�"a�ӯ���#V�x�rA����zA�{�Ry��%�����wwc�]\M�
� rB&ۈ~c�-B��K!!��N�(���D�����c��ZA%D9r�[s��.�*bꨦ���X����o�T�Q���?�`�V�Ok2��n+P%������}�V�Uc��#t��[��н^f�A'̘2�;y�.:	�"�3z0���iä�h9"� �Gׯ�)zV���.�8�&�'���P�R��vAo�1y,.�²�����g}3S�d�s�u����E�[+�V���}���7�ه	�2�1�LuKg�Ct��_���(�"=�.��]�1 �X�`w-w���eZAڵau�1�ͳm���a�_|��F�D��{�M��L8㋋���r�9�8�[?�_�R9��kKl����לB�5�Aͭ�կO�4$�]��.jr�Ѹ���~��֫�Em�X�(�T�k��6��?�a���N��J��y,�"U�Ϝ�]��6�D�����`��eЫ��)`'��z�q���[eI��������I0��P,�Z�0��y���q1�D��Yf3�l"���Q(C���SJ��&ω}�-ɸ��ɇ����:tX]<U����ER��ώ��=�`�[�%��z0�����Me.2�s2|Q�VI	�fk�׹>a������),�{�J�vH�a��E�%p!��_˽{Ʒ5����X��*[b�f��Q��3K�kXX�}�� *��9��K<=*)_��!���C�^ �@Җv 8R��D(W�8k9��K�}8�HTk�7��P��^�����7\��>ґ���Ԕ��C>	���q��}��pX�#No�����������W<��u��K0rw`�A/�T�O��,$ ��:�mՈ�g�݇��������x���*2�,�r}i�F���+��g��� �/��\^󔠣��삐b{�g��O���.�� ��|��ѷ��׺JEn�+��H�_!���ӑ��I��#�!�Uf%hL2�d���Ӊ���]8���rˇ�E�h�Z��C����'�n��������4TU���tf�} ϻ�W��7&��r��� u�%��h�#��-ӿ*@ �W<EJG����½R���䣂r�v���2�fLa�D��<����[�r�N,���o�n�+K*�7\�m�<���bL*���bMp!�k���%���G��B�����a/jpY�	�{��2N�e
í9�n,���C�O�q7� l��6o�2�ͨ:Eg���	�E:.�v�+%(`�C��{3���\����I����+[х9���1�8S���&�/���BX'�E��X�g��IIF��tZX-!�G�Oܥ!���,(�x��kN7*���y�bVSI]�-Ax��oU�a��3a!1!��	�v�+������u��,�j���aAd?7�&!�Yy��y0�}�e9}�����F�/>��	�&d�	կ)�C��+g�~��ՠ�Lg��H�
.�y�������e���=�����?_(J�������x�\�c���2��U+:�:�IoN���?���Bȭ�������e�!x�xtG���$��2p��/����������jv��
�77�
��Ðњ�"d��S��z���z-� _��qyGuZ!��!��O�W���{ۺ,=�h&P���L�&ѻVۙǾő_��/�i��B���qf	���4�P����<d�͸K|���U��}�e��~r�/��&]7O�{��{��r2�|�(�$M����Lqd�qi��݋>4^��- ��I�os�k���|-��圐��0��.��ǐUV �����J!��gB 5�S�GJ�.����� �����{k"��I	z�A�^cy[�6�Ӻ�Ph!6{~����w��Yy{����h&�jW������<-f��\";��^��SL�+�y�ctoź>�����r!�C�X�!�_G|;��~+�.ʩ�����y��;OzH�1~|�+|�@�$�/���O'��jc�`sJ�\�m6"�J};�XН�U��ͬ�|P��j�I�n�>���[�
%��%��oy_ 'L�f	�]���6d5����e��ݹ�z�IM҆��~�3�U��w�$*�u�҈J<ꄸ�(�+�'�����Y)��~]Yzs0|��G�Gx�Y�%Q��!ut�^��R�߳��=��]��TW�O���"��Sy�ڈ�z�-�u!M�ʼ`~1+\g���~��ˡ&�fô0��4P�R�y�5�`Q�ۆ����L;�-����s	����y�./e�������_u+m*����ۣ�%��8�5�4棫���]�y�n@���n�w�*]��Y�����2|���<��GR$�Lp�|q��x�b�eeԒ�gZ4��ܸ�E6�c�/l�I|,�6�5����#�{E�=Y�\|Q�GBs��F�lx�&}1eϤ#r����iڈ��$yx?��g���;�]=Y|O�:��2~#�na�V��;���s�1�g%�I˜�W-S�T�1k��)v�_K�����^�f�.		�ü�_ݮ�AC6xԒTP
�?�4�VWUs|����
���F�;�}̀�$K=\߭��D�����rC+���	P�B��#pF��[ϲ���s���7߬���`�j�T(�]�I"nu��XQy�0(�)7��?uͭ8� ��#Ól��x���d�I�CqH�<E��}F#����9	���S�h�:WG�!�Ĭ˄JN �:��~��M����d��g�&�����n��g3�3*�Pp�]*&�p]�l(�}���1܂���}驦"�b1�7�$�/PhN���U���\2�|ؚKǼ��%�ja�x"�?Fg������}%��n����5{rH��DG���1;�.+��ȫUD~ �:�$i��d������fk�4"ᳰ�('�B���-�u�ECݣ%jg(��qX�Umo�s�ӫ�xn�4� =�r�ŋ�kJi3�!aE范���V;���jA�����Z$�6�yá��.�xiwP�4��vRM����{R�B�
~&*W-�w!K�ڃ*�W�4����!��nOcZV"A@��9��
[NX�.k~�C�B����$\�o`:�Q(2���`s��O�}ʭ	ޣ%��Y�"�c�?V��4��#O��[�4���{��<���";4��U|��`-3�S(��L�c���{-[G�6�)��ۼ!P'8vw'o��"���͟ч��스.�-�t����c�3�2��0ը�:P���N�
�q-��T5(����
���og�Gr:g�f̛�
�F�1���th�i\]Cfg�S��w�>��~�uK����~���Le4m��:�\g|	�@��,>ɖx���v�f3Ͷ*�Hr��T�3.�?A�g��ن��lI��5�����5l�����;OG}5�/��I5��L�«w|��eE��X�T ߟ��ˀ���#��ݻ)���H��Jwiy'���q�W��?Di���R�M�R��2�㳽'��z�f~�&aBeĎs��o��ɋ��~0��),?�^��y�<�q�5f����fn~N"XoQ#c��&s>��1G����n^��c#���t��k�]7@C���$RdW��g�=DQ�[e%���+�!N~Hf��s휑Q5�NI�fkǂ�>���@�9)'Rǥ<+�a-7^��%�p� 6_Q)۽��5�;D׳YE*��f��o��P3�K�k�"�ͺ ���@nܔ�-K���)z��!dxC�
��gJ�1��34D�,fTWe�9������H/�a7��_���=������>�`{�[��s�CyF�[�'������ϊ#	��Ǿ��K������Ū*�p�Fsnw���/���o���8u/ j?u5�m��r�b���ywTڑo�ꄽ��*S�5Bg/�}Ȣ�{�Ќ
$��"���;;��oNJ�U%i�+�baOR9�A���|�=���/�E	��ַ_h^��[4a���~��I@��'��\urU��:hGlidQ��D+6�x?��3�g�b:Ҟ���Z4������'�Nߺ�J���TА����5����j��R_J7_��-����Pu;{7�C���Z��-ng@^n<�D1�n�>�ݺ��3pv�]"�v�vW2Ey=a��������<����lm,(�J�f����8m�m�^��bie��	M�W$k� 9�`x�/0|�>��@���hcaJ(ZY;��{`��NWs�
^�9�5��F�h����qR��8l�o
�C��Eb{�d��:�Tv-I�%�w:C�{ne����6�ڦ��U�O[�X)9��1Kq�SkF�&�B�~�|"���� gX�jI�?��
X~YG�Gn������sʶ�!eNR �br�\j-S��ȫ0��-ļ	x3J^<9�	c�+~���*/����e߇��J?�z�!􄫴_,�0s��R�}=R��󆗊���K�&�V�*����+�ˍ�����kM�+�f������W�z�֠�Ւ�͇���f_�s��=K�Л,����0�m�Uƻ��5�Lo� X¾-��ȭ�X���#E��#e��x���t�2�㷏��M2�����ۻ6D��j����7R���=�ѵ��dW,2�`�n�C//-WÞ�ᇱG�/\��2��𭔅�t������k�=k�`P�lHL!'M�י�AC�����~��d?BR#qa�k)Gk�����X<��K����!1�� �}�xE�6nr�
�5<E]���{�픳+�l\�(�_$�{�s�oq��i�M��z^2W��`OI�| �����;,��\-o���n)d`�ݐ$UQ���5�XJ�}C��\�5���SzTËi=h�T�� �i��6�k�׳I$�AR�cT�6Ȇ+�낓!1��wkr�Y�ki��kh��W�Sµ9~�-���t-."���^צ���V+e��c���U/0��"�ͤfCOG !�ܲ��H;���f�C�D�������/O5�c1��UĦP�@��/�8�����炙LI��G64�<�"�XF;�BD�^NF�#�l����z���`��n������Ƣ���� �:oԎ$'��	�ς�Nͱ?����e��ݴ�z
�L�A.��s��U��R��S5�uo�`�EG�n�J9��B��A0��4�=��s�z����;GӘ@����T�t�������=d'|��m;Wa�"�s@Q�rp���c�U�d�<:M�~�`yX@\B���x� ���\Ï�k�o��R���0�>ڂ���7����IL�_ZȜy����1-!�t�p/�Z������zTmm����`+$���%���8��(4y�7�f���'�y	|*���n-�=*���Y� ���䠯������l$v��Ww�k���xXe`�'�YZ�7l��X�E��csB��������ɟ8,�{ �zY��[Qy6s]��F��>y�1`�P��V򇞐wi)P��=^"xIeg0u�����=T��ߕ�29M�n|���;��#s�������D����&S�	�1��r)�s
KН��`���^	%�q�_��mA^m��"(P�#?Vly���0PS�i�
��%F	(���1��IKx��;G��7 ��M+L�	k��q�K#K?���������ME˔7��h����F(�����u����S�����n���"��(���C#�d߅|�E���Д�
��g��W^���Z�͂/�t��+���c��Wt���=��eW��* ��5﹁�M�dI�_P�g4�F��:�å`��'8��bw]�_�pXa^l��!۷�<�Lk[��.�X��Zb�-���/��z���,q�\����u����Ϫ%�z��s%�?���|���5"}��M�I���!��5�=HĘ�Dj�ڳyj�Ie� hX���~H�:u
ri�a��I.���1����4���`�؟=k���~gu���8�@j"w&��~�U�Xas�!���o�# 8wYO�CEiN�ha����`�V>z4&�A����0���seyޝ��b�S��w���Փ�M�t�ֶ$B���~A�-8B�K�4��e)u�����D��O�c�A[�Q9h�[)6.<����U��o��o@�QC�:��m`N!O��(����%� �}�}V����N�#*̷[��8���7��N3�;�&p�Wa3��B����^���hcGM�
)�2༜��8Q�$'?�����@L�,�M��.�t�������3��ٕ����Ì��UH��[��#����R	�O��hY�B��g5#���?% ���K\����]޺F�NpXw�%��9��u�W0����q��m"z��W�*|d�z뺊�ɱ�������A�.�el�r9H�.�0?������١�<l���n����5M���G�O��ƢӢx�d ���5�R��L>E���X�0XT{rUì���ˋ�W�?�x����1J�Xy"�X0���r�&�=D������u���8]��]w'i��zu{J�A�e?����1��y,�+0�a,��b����y��q'���`f��D"��Q�4R�d\㉳��4���ح��M�p��]2K��7]DR��&�==�a�[@E��F�����C���<�s��iQP>/I�aQk�M�>�
��ۈn)"�$� �C���aHz6�;��p�v+_�Z��W�5����Eh*��Ef�G�A3�lk�^��U�O��w!��GK��)���!�N�C}֗�g�̳T.6П��`W �9��'�s'�H
97c���qW�
������2>P���Y�N@%C�����u����&gl#�T��2���`�;�J���4��A�&wJ�/��.�c���� E�����mKj4�]���d��L�5��n����W���}���vʭ�e<^���
�6��Ѷ9 �J�Ɛ�y�ƣ��]%`O�|��k��6�|��G���/�M�E��G��F}_�̟�nn�	T3�ނ�{Kh��UPS�hBƇd��w���R���:��g��=	O��9ZϘ�����'L���u����TK�F��G��J�U��MO�7��~��0�E8u��%��m˕p^-	/�@A<�^[�)G���׾��0ԣ8��v4B'2�a�0����p���ə�tt,�ب%�ї����mwlmѾ5�Dgb��$�+��Mf��k�&q��Y��8U�Z�R��[oTaelY�,'{;o�N�_)
�tL9��סdM��R4qmN8%����oW5���^E]-t翄s:�%�vH��%�YC|>{�g{ݒb��#x��s[� �9ھz1��SF%&�)���9P�X��g�I::+�j�gX��OG`4�WJ�2ƿ�<�ߢNm���݊�7�TS�2!�c6������U3ג�W�k	�+Y���e9\�B���`����?�N"!����t0NYۋ�}زR��g������&��ե�4���Y+�Rˍ<Z����o��$\!����-��B'tN���%��s�����_޼�O����H�R�2����XUa]��0c�ou��y���P�u37��M�`�e�x���t�ё�r��h^�%�Zۖ4�Y��j��ҙ T
7��������Y|dҜ��;Zg�~�7-򥶥ܽ�G+%��{Ӱ�fM0�����0�=�P�m�L|GI��?W���ȑU���T����B�Ԫq\{����Ǫ<p��}�<Z>���,��\�?�$�}�bZ�r�a��P��]-h{r~�f�{�yi(��m$�.ƥq�7�i��)����^m	!6Z9I��I�b��d�T���`�*K�I��B��+qOUL�w����J�`�����5sTSU�l��7��e� �,�����k�E�I?��Aͅsc/�]6Z���!,w/�I�w&k�Y�{����h�m�W02X��#�-�&�ϥ"�hI^�m�+@�mc�^��?���Fl�(H�C
VZ!��.zA;rh���ߖ���{�8��O�[�1��w�!E=@w�/&�c���aܾ֧F(��6Oo���a�3Mh;8M�������x��̈́����+��d���w�FG�@~ �Oo/�H'���	�a��ɢ�$�e>�ݯ�6e�������z��u��-��`!u
ǈ@��nt����]v�ɼ����L����z�機��G.i������է%ty����=��)�=������>W�ƕ�.�#� ����j�0	L��M#Rr`t��\��ˏ�7�";�����j������R�x�+�x5��}�����L1���w I�7N�ʚ�o}./�w�h�G��S7m��;]j�Q^�%D�u8�e4�>��!"���y����ͅOnhH*�x�Y��I�C��g����O$��2���M��c�e[0���Z����E,DcNu웿x��l<���z�T�{��;YĒCQ�D�s8�rF.���1[���Z��YO�iD�e����x���gk��q�=O�*����2���n���L��;i� s5px՝" �?��Y� S]��1�U\)lc!K�|���ڜ�	�Y��yE4_SN�Ay�ZԈ\�P��?�1ҝR�KS�ghb
F~�F$j�s�]�Q�K�ܢ��x��Q�(xh+�\	��v윏#&���ѳn�-Q<��� �7U���o�`�$(�S��Οu;R#�N�Ǐ�@�.�%�ͣ��EC#9V��*���X���n�~*�r�s����c	ί�
��:^�^�
W���_���>+�@'h n2d���M,SJ�Z�gm	+�@a�Uc����q��]6��t<]`�DpS�l����r`f�g���y�3�+��<rbg�H�/���p1��G`\(}6�PE��2��%%�s�nH#?��kJ�����}#X�$2��\��5��:H��`DŁh�4�]�d՟���ԫ���~�\�:�i��E"U���3��&4>��;$�x�C�%�Cu�-����j��A���uUcbsgZ	�� o
�� 3V��?���>�ii��a;q+�aDVy�P�+cA���ߋ�여��y���j�.g�w�U��.��M�Y��1;~BW�~\g-�,/K�n������j����L����c�kAv�T9�![�.wKS�yݳ~����0o�e�Q^�/�a�`)��Otۭ?��%�d��ثH�/3VN�#�[NA���	�2� ̩c;�����m�3��H}J7�:��Ym�1�G��)����{8,y�'z��XBD����t]�b�.����j��_��3�ҕDM��������Q�8v����J�b9Zފnv�c;�=̌g���BK�@_��'P.7x��߇�]y/��Ix�w>-��������ҽq��#3���m�Y��R��|���u{���e�
vX��චO�r�f�)Je?�:�����ټ�l?��I;��M��5�N���HO�mآ�6��+�B�#�-�!�7�E>��X�d�T�%��g�������Zλ�`���TJ�`�yMf���4��Az�D_���dZ��ï��SH��'�'�Ϋz0���\�Ge�(��p��U�[�TQ0��P,��f�as)y.��q�JM��Jpf�N"��Q]��������6�����mh�A'[��I]-v����R����Aa�=:��[���+���WsK>��bsc>�Qk��Iz�(k}8�>QZ�v��)n��[��y�ac�����p��_ǫ��L�65�3K�iP+*�fjf.[���^3���k	�1��������J�!Km�@)���!Z��CX�HY�gs)X���MW�~(9 �����H�ϸ7Uշ��+<����H��F�]>#_�QL�)�sC� ���[��E���n#����AL�;��t�`���<Y�wq,�/E��HL�.f�  O��;�m�d��X[Շ/r��� ���R㻚2�K�}:sC�qㆌ�tZ����Qt��1Xc�%
H��W�at�X	�O���:��Q=|v��b"�w�E?����&_[���?�$�/����V����ӹU��mh=@dkAӺ�S��X�)g�����Zj��| �'����0�]�|�T�mЭ��. ���ӕH_�7�����1��u1�����Z��P�-��@��<V�ū��]���)���9vo-K2{��a�֌�MW�����Üc,>�� %+���t�5�m�/��xb}�h�F�oM�$Kk�l9��Z�eaF����у��a��Y1�{`8N�k
�>9�#���J�<vq�7�~1��[�	o��y֋EX�@���:_bvc�E%��CW�{�:�-r�������[P�|9�}�1A��S!
v&3W�`��?��.�g�^IU���wpX��vGP�.��M��e/�)ϕI�$N����X�	��S�u����)ȼ	;�rd�3���r	Y�+4x������ݞ��[�>�r��?hB�!*;(�U�0)���}s3����[�@U�:)�&�si� �|���+���E�	Μ�b���7��n��x�BOB���[�����_9&k
G
��̌�]<�:��㖋U���+X�o_	�4>A��'`��-J˟�>�e�8�x�XYtX�{�-�������@��q T���jG-Ù��7jS����F�dM-S���ϹE�-������G�:�6��&>؅�ţr0��k�0=�Q�P��<LׇŻ��[��V��f��J���~B��JqWg�����ev��+�<կ̸��Y���x&h}�ƺ�C�r@�
�kNZ]�$�{Me7��h^�(�(�C$^���鲿q��?i�q�ϸ^�ۈ�s�I����yW����e}t�$M�}�I���UG��뼦JRcS���5�zS0�E���9�U� ����,
kS�4IZ�XAHn�c
�76>M	�!*!'%R��u w�iYʫ��-^h�Wk0b�o�1-q��*>Q"lN^��g�+�c%�4ŋpF���ԃCń8!���Cf;Ma�ܓ��z2��������YO��1�v�ĜY�@R��/a�b� �Dט�q_���V�6jK��w���z;sw����M��"�?_����%�ߣ��l�Gۢ�Z;���o�M�'}Xq	��D����W_K5e�bhݪ���ҷ�W�3J�w�u�1�ɫ�u���;��)���I�x��7'���˾/ zD)��Z�G�Y��V����t�����d`=����^W⨪�-��;וޝ�Z��&��M�E!`o\x���Jﺩ=����e-�E�S��U�R�5Á&��Ew�8Q��$^L����R��r�^c���jzh/vs�#����r�m�ќ���Ì�%��8�-~4/;��Ԁ�
%y������n�� *.4Y�&������"7:�2��$l�(��6�����3n�eV�T�`Ze�5�-��E�'c)�T��&(�����Q{vC�Y�]3Qos�s��Fi8��h�1V�8ϵӇ.qi_��31�x�zg����>�=JY��K.�2� rn�9��x�;D=�sp?��8�q�:	��S�S��1��)�r�K�{�7��7�&	����9�_΄A�;���tP��?�?�훫FsY�
�F?����\�g�#K��ҭq����=����+�0	�?�g��#�
��<�ȳ��5���7��<Ҭ���(n�����u�K�It�A���Zڛ�H�l�둛�#tg���(��@��Z��t�����ZN��d����Ԋa�k�Y��W*��i��8G��C I�b�/��M�a��U�Ig�*����pG��V>3�Ĵ$���]�2$pN�l9(j�-8���餱~s|�����y�b�Q��q/an3�+���b��\�z��+�;�m@�%���i�j?W�5�&8��`�}�k.����ӗ#q5LBH���D OV��;�e6�o=���d~���:�5i������Eȹ��|l4�Ѱ�럳K��8u�т�Vj�t��*'Uދ�sB���5u}�ǥ .�3����X�i��a���<HV�XA\�cA����f��g�y����)�	Yw�`�ɋM�^���Bڨ~w?�-.7K�Ș��3��[����L�}�c�&QA���9^o.[�v.�����y0v�5��o���Qy���[`V�OW�ڵ�%����3�s� �V46�F#�a�[��ֽn�/�-+����;e=/�����3���k�ե��Ti��?TGÊ)�a��th8*n'�s�������-���.��L����:"3?X������Z�ˣG5����^=@���Pؚ����8)�g��~�Ҙ[�,����*K�u�]���D��w�TNʯ���)��Mk�ӝ�$���mXYF�M��|Z��0������n������RroѶ�$v?R���>��O�l�S��$�O׈�25=���9�OXj�I�ޚV���2f�6���P�E�X�RT1���"(���әM4���i)���+JH�y�~��ψ���\{D���?˯��njׅ��'�Zz���w�fe5}$�{�=��2b��0���,P@k�S�yIbLq��T�f�l")�Q�!�7�ۧ�����X�b"S�|w���](����CR�؊�\�=��c[��i�f����5v9�w�Hs�FQ�N�I�x�kXC�>M�r���)O�Ƕ�4�a~`��1y�p���_���h�5�����{�*G�2fIɉ=��3y1kD7�͋˭��E<ܥ&�K(&)�4p!�'�C3�O���q�$���=�W�+�9J��i�H��L7�g0�����M��>>�%��^���C*�H�,/ڸ������#:�s�t���D�S��8���s��7��w�.�/ b��Mۤ� �S&�m�@�SɊ���]��;���d�����
m}����l\����Sy��lO�Ѭ��� ��!W��d2�SdOccor)��l�|�yJ�=ې��K�E�oD���_y	��A��?�t�g�1����U���h8��dbD��u�8�ɳݩ������T�Z��weD'�Z����!
TApЈ��i};n��C�7p#��^�6�L	u�;��\x�Q�-?@�<��o��rS�.rK�������v�8�2q!a��4���Q�m�Ǚ��:,��l������u���m��xo�
b8<0�a�.M\��kґ�| �O��sO���"a�"Y��F{�p�N��
/�g9�JD�WQW���{q�@p�]M�6@�o�O���ES�i�u�!:�/v~�%~�C2��{����� ��}�fZ�[�,9]L1�XS��&n���OU{˯��g�ѦIp���`�%X�T�G��\�����T���e��N�>9��F�A�S5�5���jȷ'���A13M�>���	�D�+������x�h�Vlh�͢�?#V.!E�r�З�0��Q^�}�;����K����^&��.՛,��k�+S;�rQi���h�<�p��m�е��+�*Vi�Q$i��ф��_����?�! ��H-�w���1�U� ��&m=o��d��}��_��kH��z�y�VeS��x�8�t�p�����8���u�L�����j��k����7ct�nZQ�T�d�ݕ��H�� E-(�n�҉�G�oM��t��A6օC��M�Lۦ^=<��P�ϰL2���B��3��KK��w`;�Ux|B#�qRs<:�T� 
 ����<PAϸt����ee�˛}��O��r�D1��Q]#W{(����O-�8(��,$�������q�_�i��%���U^���l�uI�c����ڢ���_��)��_��%�a�nUB@|�F�}J���j95�KS;O��p�%e	 ��G�dk��IuN�A�v�c��a6y`v�9!"�P���w��SY��D�w��h���W�N�
�s-
(υ��"'��^(����+�p�c`��&���������C�Ӻ!"�-�;(zȺ��
���M�Of�1ꇓ���@-t/�6���Ғ��̘��H�.6�G���@��
};��X�/��
�}v��N!�����Zn�s�q漜��vW��O�o���'8�g	��ۜ��-Ј���etʯݥr�s��r�������1�u@��6��$�?�{�ѓ�7ɲ�f��Ժ�jv�z�f0��K"G�i�� ����tox��z��ߟ�=5�g��A�Wr\��Դ�V�F������*�a��MYY`j��\�]��!�X�ϡ�� �� �PRP�e�!G�ֳ��i�(xL'�h�-np��<c�}T�e�/�/k��2��˱cm
���� '�ǘE%z]r8��4��죗�o�%F�yzd񛃟�nޘ`*��jY�٪�����ݔ��M�m$�n���nÏ�T�ΘjeQ�8BsZ ���H��E"+�c;-�5���Gg�D%I�{1�JY�H+Q���s� F�Jid1Q����3��,�izr����&x�C�g���ŧ��=E8�ߦ�62j��n��B]6;��s�.<�ӯ;�5���=TS���1׍g)b��Ka��r��� �	�#��/N�_�mA��]�~1�Pv��?���HMA�0���
���FZN|�i"�B�K)�6�.������,�+}�G	����{#�i�G�^�c6/��V+�7�����V;�(I�C5��uqk�D��ic����Q͙h�l�#����MZ=�嬽��lj/��=��iL
�^���%:S�����T��W���J(�0Q��6�� $�1�j�KMb�T�P� g#l��w����K2���`ß+�<��]��{pIh�l����/ƹ����E����xb�ۊ�X�/������}��\�����Ǩ��%[if�d�m?�f���E'�0%}�Л�u�ҖO5��H��D{<���������"��| P~�8):F{Gi���2#� �á��4��M����[0Eu��%I�QjS#e�ݰ UY��s, �p	@@� )T�j�m�t�i���a1z��l�V����A�@$�A 6�"b0y/R��U��� w<��d}�M�����1B�);~���-�amKhB���E堷|�����`l�cF�A��R30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���<H����\F� 8�,]�(��afR)�a�sv^\�!E�׶W��ڮ�-```��t�q�8��^C��YuC|j��?�9 E~�:`r�Ķ12~Up�{��Z�z�H�	$v�J3~�qY]n��FuY�� ��.�?��7����
|���8!�-��F���+%^�X&I�wWB ���A�����
�t�-�ҤP��m�͖���x��'�Ŷ|�2�93��K�����fb�m[&�2�Nj?�Nz>��9G�:O�j�>���G_(:�^E�gT�u��G���L 9I���6؞�|!���;�tT��6����9���ܭ9���E���!�'fk��3�rw2�a�W���O��x�����n�ߡ��H��g����-�HM9��·�%�W��Y?_�-#�'��N�����b�!�Cǹ���i����l�#Ӧ0Z����.0y�b��9��mmtM�ŀ�n�o�(�i�]ȴ��I��@�cw��:J&߂�;
a#�IN�CO-���\s6w�;�	+��=��[S7a�$��c���dJ]��}����(��nG\\�p `/jcL�����D���t��<=x�~e؅p.\l��>�NE�at���;Xk����=���q��,8���ң���z��Q5/�����ė{�5$.�E���@�}��i|�2�o������/5$��ɷ�Ѷ'ѕ	�k~w���I�z��6������B�����̀�I~�'�c&{ƐN\���Rؗ[}yu+1�=�P����{�	�:��ki�w8�؍���K��j'���z62,P�
^���Jjk؞w4@v)g��rz �!�2�� ���3Dfw�e�ٌ]���8�@�d�S������܁Y���KG�ǧ1��O����#G��GB�BY����2Qv+���.P3~&,4'S��&/�q��;�a!�@>��Ik�3�K������D�'�VHN��@]&JeO��pV71����R=m{�D�L���?��`A��R����#hD������@b����NK�����yL~��Y]��e�93?ix ��J`����P�N��05/���e�	�N�n鯪���@U�K�Q)��',�gK��=yN
4�3W�`��.+�t��V�I��w�pה �"(�ƙ�
��u�����䨜3��4+:*�Q�ת�,��	�u޵�:��2G�RF�"Ofd8�NM��"gI�kҤ��z�\�o}z'mO�=TP�硶�����o)H6�/M�\Fj��9�͔/_�iH���)�yNn��0�z�4����Ć{�]���
�f1����D��B5�T���G�Ump����P>FOeL�5ѬעSm�.�vj)�*K9���{�p��$����J�f�wǶ8Q�j������||W����Eċ����ط���vX�	��HQV��'�RJ{�ĭ[�ii.{V�!�5�4E���4đTEv��L7c�����>k���l�Gs!�H��0��O��
xէ2g��kcc���, ����|�w�Ev���!�?xk�g���W
�*i�\�Ҽ!��9��E��f
��=�_�[*B��]��w��s7�-��L	��O-,{�M�c/FSG$*qa3�!W��a����j,����-0}�C\�!����������>\:��?��J�K��B�� �҆Ts]k�:�Q�Q��\��| �����ӄ��X"q%ɻ��S	��Z��c����{nZX6r����*�.:�h����
�rߧn)�	~�㸇ꁫ$:�ӟS.L�پ�a��ږ��=�(#������Wb��a�T�"�M��~�9b�
&�']��K%0O�+=aO�>�3o����';m-�<�7�������ɍ o/��(H�N��}�;����9�Tw6LL6{&�VE�H�^�mF���o*79�L��3��������y���=��l�K�p��ʢSJ�󃴇��S��P��B���hw�HSA$���YHɝ�)�92f���W�^N�6E�mn�^Vw��D���_[����T}H����)�=�TV;y$�h��8���ɰ��Qtr��8�(��O�����}��ʾ8i&�iբQ�BY�ȡ�T
�����)}QA�B���Oh�2N��W�ت��
o�o����a�քd�E9��_jW"��\p���z�2[11��2�>�d�w�	�2��3R�<���M�_1
}vS��ςDx9�>����ģi�?��]���KY�X
������	]�6��c�kZ�&��I�=o�����	nzfrj�S���� ��c�/
���$��^ܱ@��rZ��׫'��C�#9�7̘����ݿK����5���PÈݙh�dZ^�B��q��b^��{={Ep&O���:����ޅ��k�-�Es	v�t��&��sʻ�8g[[W��<�zY�!��ysj����Ŗzz�ա?M�
�ͷR��(ե��r|ԋqd8|�-kٻ�-M\^ �$g�{��b'H����_��?��w�y=��b4�
�U���'�	6,���y�;��Ágv�-�L�4JFgٓlH�j%�)������b �/8F(}6ӌH�R�.��r&ܰQ����s�8�Dr�>�S�Q���q�ۻ�7`:>%-�+��|n��4�?"��W�2Xi�z��:���Ba��#l�;�	�zC��� <�E�5�1��F�/B!hX�L�]T=��M��G厽�s�������0 4�i�Ҽ*C�_���|A��.\h�HHT��w�W�*i�ܮ�:ׂ;�䣺�V�CLX7D��*����� h�B.'9ilP������C}2��(ߵ���7T�����^"�]P��Eut-��^A�"<����|�r'a����%k��I���Sfx)9����E3��B��[ �G�%
�k�g��i��Ia�V?��> ��w��J�̜���\zu��;^�	��΢�ѿs��H;���j"�21���-�-{�^�W�C��IpOlF��ʉ�PE�YJLʫ�L?0�?!��V�Np�a�F�t�%�&�� ��JxK���S��1΅��JH\�W�'V�U~_�3�2	���w��G$�	�"��l����f^�_Q�|d�I	����dq�9>Ħ�稇l =�:����u��ȟƫ	o'�X9��~�q��͖��a�O��'�Ư�����!�|�&�}Sn x��^u�P���U�yed�$W���vB�.7�\ 6,&E��6,��(z�D[�4)�I{���ܿ��>�����5%tH�(z�Q߅Y����r+��>ԕ���2��Ǫs���<|X%؍�bb���d+y�Z�f��aEC�.�F��P���f��:s�Z_�^��{x6�|jb�.�&�<^K@L}_ȣ��C)��{a�# ����o����y=U��iv&��� �in0�ay�u�T��MCU$O'��&�B%/ȣ��'%���G�U���5����N<��]o�/t��4�o����S�U*<	I���La�<�+�鞃΁���!�疒Ѷ��`�	���N�i��̺Zk:�����0ͥ�f�{<��'B�ǂ[W���ב?��C]hB�5����=���9��d�+F@��do��Z0�J�a�+���3��t���-#�����h��^�LJ:���m�\�D��)�����`������E�c��2��(�(q�,�2�(���I~�l6���p1���'_Pl+qumĶ&yJCY�_��#�K�hLg��ik��5��	/��X����;��K����`���M�\ݫ%W��f��X�;}�%��=�Ia�����^%J�L����*d]���)�M�LD
��D~�@?��|�c���F-8..�Vl:TQ�v���X�q��������4h~}.C�f9Ͽ�H��z�/ٿ&�X��*��ֳ�!����f�I�K��xx�Z[�G�<�uТa<�55�8�8�2}������,�Π���ӆ	�N�2R��P��S�	�<���̍R��?_��^���g[誡�!N�Go�,�~�^%Lts����B�gp�l���������A�����tEڶ��6���\ +�4Re/��A�"B���~�� �0�~]g$j[��%���:q��^�Q/�(�?�T��V��5*m�7,.��ql6�A�(�
M{�`�@ <��5����c/oK�4��֯v�	�ƨ�����Py^R�����O�����3!�܂}7���/��YL�6��!m�`w%����ajV���<�
�ۑTn��M�<�6�������՛��s�{�j��T!��"���m6�S�޿H�؁g��2���a1	t��Hl\R��8Ī��y]'=s��>�v��A"j�8�5����I˿�]�e "!}/�G{.-Z7<r������0O�^F�-^؛S�YD)oe-�\7��<]���`����p����pP�D����/�>ֈ��	9��{�3���+�TV� ���XWb9L����젊���U���m?��M�϶����>�-u�����p:.z=����l��L-��3���#C$����e�ڜ�Rs^�3�����8O�۱.��˖!]���'� fv�RC���_�d#|���3���	5 �\MR��U���:�0�gy�%:�<ެ{S�Q��>�D>��|�k�g�Ay��2���K�K_�喾SڙgT2c���n�����7&O`s
�9TS�؈iܥ��/dZ��-�*n
��`q8'����>�Q�>�v|�0h�-]�������X��M��$鈄�.�	<s̈�k)3Qpn5V�D69��jY������6���æ��(�ަ����vOn�d�ϲQ��%�q&�@��僸2�>�����h�n���S�����;��1*Ȋ�Fi�a!��y@G���S��R����ּ���pr���Z�����z>"���Rk�JZ��g,;fZ�o�Ҽ��_"��|�ѓ4^4~ӊ��| L�-UoF&tps���� �גI���
`lJ|zo�!ͻ)�['�ԩ�֭
t7K��I����7����Y���#��N$$�*��*���߭�R0��0nQ�:��#����u~2u�sH4����\�9>��0�q�U�
��o�~!�0Ɗ�pbka���Jª�"�^�HΞ��׳�^X�A�U���	N���;}���_�Y?֛�8B�V})�j�h��)�!�1r:�s�M��^�vnaqU�c>I�U�S$��%��>˃�D�����&Cc���>E�#�\{PP!�o�ǘ	>�9\��W����D���ReBL�q1q���½�*ɨ��T��� ���!��euCo*%P7&6S3�?�Í��N�NW�5Y���1�L�m�r#?bE�D�N^��J��Iu-�D�ڄ9L9��eeJ�8]��z�Tߓ�&fwH^,�O�j��E�)�� �Y�8a��P��������AN q��sn�� ��x"�1E��)�)�͗�t[� A'%������JK�Z���;R��Ͳ�y����]���w�s��F�(^x�Z<�3�ʿ�l~������.@��碶��v��s�}�DH�8J%�����B?�:�@��YZo5F��%�uO�Mo�d��[r���eS�����[���\�^����� � �c�?e��hH>j	8d�[Rb2�	w�dl��`5]TNv�<!h�Pt�������Y��������%5`��ij��sh��L�����W=�'SEv�s���q�=d�J��aH��@��I~e�i����������ԍ��v��}�~C����.�뭻b�1: /��b9�ĝvo�H[a�R���k�_�ZЏ��qlݮ��H��n��Լ���F5��u���������bu@l��#j*���o$�}��b4�o�3nXwY��j�r*�l��Kfa<VTۦ�T���ȥP=�w~^]|P�ɻ��g�Q7��n��Z)��T��<�P�S7?�*Q�䗖cԌ#2���A+��r,v�޲�������%8G���z�+E3���j}�<�<U�8�F��8��b]GQ�ʎ�g)ΆђΆ�s����T�n��ףw�ք@��Zw�`����)����'��?�C�$�,�z����gT�f>1�19p�9չ��Rz����ů���~%C�];|aF�)g��T�ۛ�Ut$�q%y
	��e�^��AFf��+2�}X�Ew���n��A%�L����~���]U�mM'��mx�����C�2�f�����Q��swhmݢ2��?�d�>i�G�J�7֢�I)_��Ctr��[�-Tg�uy��G��+L����ثW�!bs��<"T�D���96�f��ũ�����.~!�|of�kW� 	r����\��PK��,�����p����@�������*��e|M�K�֔.��U�m�,�C-�������[zbE��C�<#�uN��3zx��M������9j0F̹b%��ԭ�tɎ�^<Լ[�1ݵx��d���Rk�՛@�`�����JsS˼�8aa���Nq]-�h�ɟ�w�� ��&kΊZ�[@ҙڱ�Ic(�]d�#����V(~&�G���pF��d�cyo�註��!W�t��=�-~�C�p1O���-{	�aAaʨ�X���|=S�=�`�ڞ��N��DM��A��p��/�|(܎4�{К:$dEb��ľJ��i飋�|�u�L�
�͑l$�B*�D�j�9���֝�~�~�V�w�K:�6����� �B.��1n�M�9~ �c3`����/�� �؄AMy���j&�P�P@��f��-O{�đ��zA����+jT�k�GnW2|]�i����j�.�w!,�v��k�A� ��2,$����D�-�PC�J���~��mzۄ %Cь�m���Yj��������1I���dX�����oKGO}YQWK���+ϔH��3���4�~����į��lnnޱ@l����|F3̎A�U�k�h��D�7sZ�NG��@JWne��1ҝv+1����{�6^�#�"����.��Zޅ���h+�W��M��i�'K������k�7�f�r9�X�xA*���H��b�;Ι�:��̸veæ�Nk���������3)�>�wjE���Ȝ
/�Nw��3dӇ`FfHx˨ØI=��H
 T�K�3
��% uH���9a�������:W������s���Du�R�:� �G G�Fo�O������V�1^gV��|��B�\��$}^�O��T�'�#���7�)�]�|y�\3 ���R�=i�a���,0�$>)�-.n4@��m:zC��������̛$.`�,��%�4���"L������rUo����Y���i���9�5^�>������Rj�ӆKF�i�(�ɢGE���{��� �8��j�L)��IK|�z��E�x���s�T�	6�CT�	FH^:|�b��R��Ě�5i��V5n5p��������'��6dZcmm��k���l�=��eNUt0Q%HOݣ�x�E��Z�k�0��3��m|�њE#3ˆn�9xX���j�
�Qi�L�)"�F�kE6�
�&�7����&#~���J�y��7�*��^0���,h��MPv$s��$��qz�4�.�:�?n�!�8,r��Ѻ�p�������C(� 9�Ʃ�>�?��,[$J,�%��`���ۂ���	k�E<��*��7_f�il��Vӱ�X�Ѡ%66��`���#���z��d�^�r#b���z�:- d�b쭳0�r,�"P=~L']�7��v�:e���3L_]l��m�ǹ���O��L���`��M��o�@a�53"D���>9�r�&2�jݱ?�O��a�U���r�3\ꖲH
�;�y<�	9�d���C5 ʣ�H�H�錵v;C�x�������LYl��aVc2�H��^m�6ڜ0�9����R�����q�������m� ���x��py�s��nأ��4E�S1�����)Y�o�ޖ�VkA�����h�J�W��V�p^D���Ȏc�m;V�(�Q
Cɡ��ޜ���^�������
g�Vx�;�h�� �<̊�z�Q�D��(�Ԋ������B�}3��DS�VL��/4�B�ൡ���
�����O�}��(BѠ9OU�3Ne�%WJ��w��
�Io�qz�q�#Zd�Ŀ����WO�\=�t�D9��?6M1x$��`d��$	�c���a�	��[�Z(x1���v�^�YH��N�=O���������v?�ЦT���P �>���Q��z��](�O�����1&�o6�=�k.���	;"zr׏�S��.��S7�K*��%��N���@��frǝo׸�[�/Q�#�K̅���!���x�ē��h�4P��H�29Z��g�/~�q,�5^�=Hd#&�f���0�<�x��W�k�x��=^�s6L�t�/-&���~�8�WW��g]h!:g|s��4������F��!�Mn���oE����8W��d�q1�cښ����j3M	=�6;LTș>�H'=�3�Ĺ��ri5?����T���X4l4���U.��'T�,Z3�y����8v#y�e��47�� ��ƗLH���ǎY���'2%NFu(�y]6R�w۟*J�}ۗ�R¾s�i����B��7�>O������`E�-O��j�3������D0��Yz�xRٗiB���p�xfҟ$��{M��`)�3�)�ܾ��|`"�5���*�!��z`3yF����j�l�x4��c�n��aM�m6�JۗEM���I�-{����" ����f�V6PcbZ*�H��Rg����p1�=y��m�{R�th�ug�]c|���e������O<"�p���Y���q�{Z�]!"ݟ/��^.�Ѭ7J5�s;��!O��[�i����D>We�cC7/X�<�>��D�ȓ��He�,k�D�Gt������o��Q➷���$ag-�VL7��2G|b�{��f��\��惊���6�8�r����b��&��5{�p�>�= D����ňTn�BA�
��.�?-�閩�R�3|�9�ܛ�����u͖���	 "2Rڭ�l�ad_�X���-x����j����Z����0d�ay%i:�?����hQ��v>D�.��gFaTy,����K�!�ʡ4�S�1T�.xG~��*���O�7� �`�`&~��SW���Db��;�bd�2-�bnƶ�`���\9��H��Q��ͺ�]��{-�p���'�[��Aߣ����@��j�g�KX���'k���6�5ecr~���cY�������r�������觹�e���H�28�n�dL�nY��a�7&�'0�!B�2�Zٻ��ڼ�M>n�w3S;Қ�@������͑i��ӻ��{@���Kd��c�#��xbQȬ(��H��Z�*`�sW�"&l�M���~'Z\�gC^�f��o�"��d{"�u���z4�#��FkL|\���΢�o�s�t,H��tM U�qI0\�
?�|���!�-�	��zV����7��I����t�GӚJ�#���$��+���ʻ���it�ow0N�;����#�L��1G�u�S�4w�Q���[>���0�U�p�«��!����	��k˗�㥼�f�IϚ�G�Z����k�X�FC����������;9v�c��3��t*$�֡)ʾ�hulp�]!Tr�����_!���Ev���U_�>��P��r����������GʋbP�����>�cu#�0P�l&o|�i�EHz9ۭˋ[�l�H�-��O�we~>�-���\P�qYT*���C��\���ݓ�e��/*�7b�6}/?1E��;H���ƚWn����1����LK�m��]?�B@Di�@��%�9L���@��Lu�H�!�\޻�����#���q���.u^�_�O�Ej��k�[���F�t����E���ז�2 ��d�/���<% x�)E	������:�0�1 K��%��	�����^Z ;H:������;���,�3#>���(	�Zx���opl��Dn2K�j��գЄ�7\J�/@���l8���B�u��|��Y�CF=�|%L���Dop끗xƊ�rS?��ҏ��[�Ͷ\S�����ܼ� �~�?!.Uh��	��[����\�ȭT��lP[5��v��|h
�?�Z�,���Yml��S `���l5��(�%�?A�Ȍ�Lv�h)H�x'݊�O��s�#���q= �A!f\<a���v��酉V�%0�r^�z.%�.$��j~+v�qq�����=�.�Zu����:�<7Þ���Y/�v��n[$9�$�#�g��pVq(�,�OC�HK
�z�x�B���jބ���9�r�v��b����C��*��C����Lb�U�oX:Nn�Y�w����&Il*� ��5<U͸�bLH���'�;0w�c|���AW��Qst��_B��ι)O��3����R�]?��Q�S�+~#n�	��7�+�PS,������v���v��'p8�>K��k�+�\T��I�};��<!ti,F���8�,]?���E)���
ks?)XGȈ�*.�����@*�ߖ��`U�����o*,�ʞwC�L��h�i�	ߣ�n�"�E1��p�����x�z���2`~���B~a\a]��F�0��"I�������;l
Ņi��dp��U�F��[+�T�Xw`.��!�A᳒�"�x�������m�vj������!���O2T/�@����ܢ�/�mD�2�y?��`>%��G�^��8��\d_HJ������$THm�u5s	G�PcL��ř.�E�g�p!�6[�Dg�T��B�G�梒��e���YN�rv�!ͻ\ft���\Era�[��٪�p����~^���Toߪ��B���e_]�3�4����M�<��B��s̋�h|�-lf�MZ%�fxFb���C�xiձĚ�<�>Y��yU���*W0�Dba�ǐ�t�Su�����q̹�����g���@����MJ/f��1�]alf
NTZ-Dy>��w�%e��M5�Fi�[|���m�WcdP!dӹSYk��~3�(��Ge՗pI�hZ�c�Ps�d�յ]wTtz7Y=MV~nJ(pW]�HW��f�a�+��wc�`��=�t`zcg�>��;���B�ʬ	/I�\��K�{���$W�~Eye @�:i%8_�8��^����$ٔ�� ���uSh����~ �����I�6������B���mh��	�~\�-c�sې7������}y�`7˦�NP�A%I����u|�iV�怀ض���[�j����[�2��P�uu�ܠOjt<w]n�vr��� o��2h$-�q�D ��n7���Ke�:��%��	���k<I�?Y�Tz���;�1���P�s�C�G�Y�N�;}+K��րV3���4�[���Ht�Ͽ��$�s*�e@����[3@��ƅ��`D�/�?I�N�@��eQ�٣;1z�%����{Q�&���V��Y.�Po�-y/h��&���1�	�g���)K����%���L���\��"R�9ܼ�x�,��3�k�����w8W�y�6�Z�eorN����s�o���^�E�zl�3Ю���^���FN��P3 �e`���4ư����I�o���� z��o����u�����K�Ũ��}:�ə`{a�g�q Quǥ�:���G<Y+F+UO� mЛ�/xg�p�mK���.\5P�}óvOL�xT�i��_����)1�_�8,]\o*.^���y�,�k7���L�a)���n��B�Y�fz�2�*��M;��
���E�O\�箺��6��liu~u	U�K�|�=�9k�X/�u�M5�������tj��Kg��d���華�S���*���X8�2tj:&ϊ	�|@a��]�Ĵ:��/���E+c����	S7�H������RS0��ֱLi�I�V[�
5,F��1T���=�g���Zc���;Ik�lC�`ʑ�(q0�P\O�6\x�/����k̙�\0��Vb\|��^E_��*��x�_�&�h
V�Di}�Q�e/c�y�Er,
�{��<�)5b����m�ҵ�"7s�m�5��X�~,��'M�-��$���q��N�ꋘ�{/���{�,�n��v�����i����9���L���A�>e���h��J���,6ԩX�����k�ၘ:>���ف�>��Dp���X�J3%r�b�i1���4�ln��#�l�t�r_/0ѳ�:i s�	��;tr��R=~9V�S����k:�S��$�L��A�jL�� T�X]܇������ى�;+m&a�8�"خ�� {9�|�&n8	�����?Ouo:a8ճ�G�&3�(ȲC;�6{<�n�c���� X���D�H��H�g;��idō�8L����V�?H#,]m�����"9Zu���Fz�S���fڂY;�9�l�܋x�-`p5An���a���p�S�����Ґ�ы��c�A��r��9FɆ��Bi_��x�O{q��gm�S�V �^�zF��2A��_�7�#� 
��8 �Ƴ/V��Q;Bw~h�����DQ�����(�����´}��}o c�A�ϰ�j���rB�}{�p
a
�~X룳p}:��B���O�{�N!�FW�,��3�
��1o�-e�ѻߘhd�Q�A��W�Yt\����������1����K"d�%�	d=t�@����y�����K1���v\��GgW��$�y��}�x�7O��2�_����<+����s�Z�6�]d�VD`�T�>&��%r=�9+��X	�N�rT�Sd3�ƪU��Xr��{+��q@��r�j�t���k�d#Brl������U������O�4���P�f�Q��Zg���k��q�b�^R�=��&�K�!D�x��ގvek�n����sr�7t�L8&+Xm��8P3�W�q*���N!� 1sӶ��D��?�S��YEM��Ǝօ���������јq��(��f����ME���M��25�XQ'y�R��ʮڮ��?�$�ܨ�C:4��XU�z'N��,@Jy7iX��d�_�!�4s V�܋��-*����Bys�v��nDvF1/7ӵ;�Rֆ��ۇ��9ࠎ�^�sc��-`D�G:F�z�㉺5a�$d��t�o{[�Q��KI4��%d��_-�� z�?�/bz� C�o�����H�ʧ���1R��yn0�
FbZ�2ǩ�t>�)s�׼���
1`�ɑ�xV��K�@���z=J������aT4N��-1��z�w�7��+��Οe�[�? �~c�d�:�Re��N�(�G�G��pF�"cnC��=p�V�7t�[�==�.~��p�h���߁p�a�$z��唫y�9=�D��:F������b��Y�ʥ`[/bҿ�E�{��$��E�8�fߕix��QP���|���$R)�ə���.��k�~��+b����6��Ä�B�Q��&����	d~U�c� �p�����f�9�yW���_��P\A�B���ϩ������ �/�D�-�jI����#H2��"�؃�g*jͦow֦*vV��=v HQF2a�;��z�D9����<��쓭��b����d���!ab.�Y� 7��#�iF�1�p��7�)ע���G$�XYƏ����`+��C�oc13��34�H����O��FB�]JQ�j�@!���+bX3����S�����D���x��N\�@�J�e��Ғ+�1SrL���{j�����7�IߍCޯ���)h�Cg��/{�"~٬�h�KY2���S`S��{6��b�9��7x�ת�l�ۂ�c���4s��ܟeXIN����K,�;4�� ��U���i��(}���*N��39t�`�!2�-�xHIpQ���� ��m�h����u�NO�N�A�>d��IB:L�Q�9�������u X3:��G�}3F�O�G�t�!(�g+}o�H%��;D\�ݡ}\��Os�T�0��XmB���)j��ꑷ�\� ���6�2 ����I��_e�W)!"nI�[��R�z��Z�ڀ&�����b���Ȉ��؜@��$D��?ʈW�
U��#���r������Z5�}��uZ��}�j�U�Kl�ݝfT�\�ٯL�ҮH�����(8��Gj34pϣo|y2V��->���`����|��m	LOGH3����^R�qB�O�iKE8V5�_�2'���v���K��c"Um��͍k��l���{�*Q�0ƜO�	xwn|I�k�Z��5��O5|��E�O����xם�E�
$iVz��^�޳��E���
�TT*�=I�1�a�lҮ:37���nŶ��G,d�M�DhPm$o�q�.Ͱ����ں6s&,'Q ��"�e[C���$�2S��ea�;Z�>�������J�mN��C�ԂC��D�k�@�s�A�Lc���ݳ�Ӧ�2X��%kA�5�ح-���@�����<A�r�	ьF�:b>��g��(��rA2ˠ7~��������:�no��ULԡ��ð9�|�E��;�A1��u��ق�D��az"1\ƔnY�9D�`&'�Cr�+��{O���aq䞦��s3곲� �;�:]<Y����[ ��0��H6-m��0;8Ĭ�B�=��ָL.�I3�PVxxH���m(wڑ;93�|����l&Ik���*�粬j�u6�m,�p���o����g�SF1��K�����3Q��pA�e6���xɿwm���$�%����X\�mл�V\��&<I�8�����T*'b��2}���+V���;[BJh�X�Q尽�\QV���9S�(q���+j��~%}�w����"�t�ՄR�B{��I�m
���뼐�}sB�j�O
�&N��zW?!����
�ޭo�b�j�8i7d������YWD��\�<��y����<1�ɢ�uddMj�	�B��VJ՞
���B/x�1,�5v����R�&�
2�0V�R�0ԣK�N�D����E�AϹ:տ���Ɯ]]��oN��B�&-���=Q����&	��wr�FS}F,�@��`����nsٿ��@{T�r�Z�׍a��/J#���:2��v�	�mp�(l��P�:�����Z�����q�lz^#�=�X�&�����O噱����
k?�"꒮�s+�t|��&$����&8�M�WӪ�\�!�<Os�Eb�T��8�ӄ���M��Ҏ/0:�:������	q�M��pŻ��{M~T$KA�	�U��}'2�Yڧ�`?�vi��q^�m�4Z��U�[�'Cz,� �y0Eḥ���M�z�4�Pn�u�0ƌ`��F��;>��b��+9F��V�.��RoO۔c��3B���s|�-�fp���Q���W�S�U���1`�ag-���o ǵ�4}��&,��q�:cz����,K`B�?#NC�+�z�쇰25�']Q�S(S���B����.ѵT_6�o��y9��q���%ʘ�35x ��i�`*�X��c�:A�͏.~�O�s��& W�P
i����t;�}׺�=Cn��D,0�Z&aۼN~�L'��MP;���U=C�}Ȋ�{�?��T�"�ޛ�^�tPP)|�uV^��O�A䪦�<�^l�Io��o�;�ǉx�+�����xf\�N`�'�@�d�[b��d%�������xI��>�����Q�?�K�����߯�u8�V^����������ƣ]+i"xk�� h��tp^�}�Cm��pq�
��и�k�Y,G1�У�0�z2�j�G�0�����G�ֹI��k���A2J��@�I����ޏb���J���WO6�V���_�#��ȝJR�w���$�0*Ä �lXW��H��_s�2d�J���ͺ�FS�9`��I�l�k,�<�����66�M��'�?�9'�`~�o�~(��&�q!Iv�u�Q�V��Y%؞���߹� �@�r�Ƙ�ƞe�=$9l�f�.��z ���E�X�#�~ ��z=z�[����o߲T�ſF�D���U�W��H3t<z�q��g����#+��7�������k��hB�޵3XF �--�b�/��i��y��f�D�E���.��Y������	X�s�QsLL�@�D{���|�sr.ud�Pq@<za_*�����)��{�$� ���w���-�U
|�˪�W{�KC��<y&M�0���/�_UAV�o{�'�;&��/9;D�A���^G��c�j���~<��$]Qx�/���4_�؁�ۯ�7$!	k�ʮ[�<�H��˹6Σԭ�"͖4�G��C	)�NF��k��ZM��3'��jY�4�{�I|����~�<0��0@��qh���5�����}�Wz�m���F۫(������Q�J��+ �˽Vw�xۯ�!E�d�Q�B}��EO�*��p�i�=ۨ"̸�v���$�_���䶟p@��X�~ʞ%������G6�=õûB��˗��s_~��c��4�aD����q�jj|y��� �P�|��ܼ��;�����`�o�~Yfj����m{c2b��Xӥ�ij�^�wa0v\V�&H� ٩D2\�[;�D*͖��F�0H��$�6ӆ7�F� �r��30JY�\f�S:��B�1��1w���1��U��G�ְY�,��� �+�[?����3��4��y�H˹�T�NH��&�@R��|f�32�2�{���N�\D��oi;6Nm@0*�e;�/���1��X���H{;�oĢ��HX|߾��� T��W�Th7���=`����@�ωK+�����/��0��go��T9�:�x�_��]|r��d��!{B�c<��2�e�NQW�]A�,��Yj�$�{�h��U�0� N]uK3
~�`�e���J��	I��h��� zH��~���u��_ƅ�o	j�g��:�Gܙ��Y��[{�u�]:#y�G�æF�O��m��1ٱ�g�I+�Z��&\���}��mOv�PTC�f�	����e)[u��}r\��H)��x�͇a���M6-)K�nZ
��|gz���T=��綰���|h�y<>��{q�űuT�EZ����@UU#'fb��cՃ��.5O̢�U!�j|�K�}�ݎ���ma��}����9_�
�8DQ�j����tjc|jߖ ���^����8�o�z�i��	�,�H�e����R�=�Āl�i�Y�V��_5����1!~�O�ghs�\��cSD��%�Wk."l�Npt���fQ0�lDO�Gx���0Ak�����v� v�|~
\E������+x>8՝�t
�e�i���M��K�E�@�
(����'�a�����G�_�37]ƣ�_���,N�xM���SK$ ,�q`�9������s��GE�,Xe��`mξ�?b� ����6q�,�>�Q7���J��S�V	�����*�k���d�ɷ]7r�OI��.Ѐ�M�XM�%X��Э���֕W���u�'r����i:fw]�l��(rR6�8�~�,ڇ}��~�:K�w���fL������(��B�b��z�.	�3��a�"B4U��3'9�&���E���O_��ab�i��(�3Be)����; F<�b��J7ӫ}� �Y|(^}HgI��2��;��6��"���oL���$��V�t�H�|fmys.�	�9�����ܯ�=ʳ�X��b��
i��; ����p�����~�~�級�SW���|>������|�Aw����ɰW䊬�w�Vw��9�����]ma:�Vʬ
���h�y������t{������0dV^a�;,�hVˇb쫰��Q�������(�����$�gg2}�zU��*�<����;�B����N�
jP4덺�}d��B�L�O;N.�W��؝(�
r��o�~ �{��I�;d�{��+PW�̘\c���*����,]1����H�d~�	N=��j�/��e�S e�1|�v�\����wn�c>�4��H���F�,��� ��湋��l���L�]@�T�~��&>X��=�&�E2�	aOr�aKSN���17�qz)�����r��A�@�Mr��4�^̄�:#�a��k�����2��7�Ĺ��N�.Pvl~�{!"Zѭn��oq�d^|�=n��&qw��x����u���kp_���!�s��`tuy&Ս�}�=8z{�W'�=�M��!�pMs�'��������{MԅÎ@�<�k���ަk��qW��ڀ���~zMoD�\/
:A�<T'�����P��X�o?w�d��ȋ~�V4��
U��o'x��,��By��Z�vw)��.z4CC�������״���%�`[��>aF�n��_huR�H���wܣ�p�8дsM4G�W��C��$����A)�N�|`-�-5�7�@{���	������*G����zH�ٽ��B��#Џ�K�z�W����x�I���R9$�Bt"	���%TP����Ҝ��PE�����_a��|S ��8i�,*�NϜ���A+�p.�7H;
���w<W���i�=y��Z�;�֊��[C�
�D������ۍ~�'��<Pl˨�ؕ�C�H�'Z��0eTi#�϶{^���PZ�u�_���z�A��V�W��/�[:�� ���Ů�|Y��U�~x��\��L'�I	�U��[sn�c�%=#�����\�eIX�߈�oG���Pʅ|�j��W��P~u�+^3�d�����&L0^ɣ�J�"�p��(��� �^O�jC>Լpb���C�#,�Y}\�A4	0z(�o�'��t-��8����3�"JB�ګ�kM&�W����.J���W�8�V��_W���%ix��w`�$�S�Õ�Pl��:����_�2#ds쁱;�����9Qfy�Z��lӯ�D�!!�Ǯ�����'�ʃ9�(~"4�c}�����lP����^%�؏�(�� K�K��H�����Hk�e��B$
&��.�] 	,E0f���R�y�z��}[�l@��wy�e͠�w���Ճ
��$1H�^zf�L�8�⌰A�+(L��h���eA �=�3����O�X�����b�7�Ԛ�>y�9fc�YE6`.:�E�b����4�+�s}���u{�|]-.&@��|@-�_;�-��ͷ)�{�@" ��b��s����U�r��5ڈ�hL�������y������� ��U2����8'ߝ&*.y/�u�ҫ �A�aG�����*�<��x]���/��4�6��R;��z�	\�|ʿi!<�z�����-��Z����z��	��NW5ۜQZ���㤨��#1���{��r�:N�������Ni�
���u!8h5�45>z��j�����~'x�w��y����/��MLJE��+�X���ӂ
�I���@��З�_�Q��J���9��\�yE���j�w���N-Η@N��Vs���(�i�q	�/2�0�y�tI�� 66�c��� ��_ѣq�hI���nC,���K�KLZ���(��_�[�o�/ ;�XaŶ�nΗKg��S�W�)�\�G�%jfDf���X�7}ű��/IT���=�p�%]� �r��ت�"�{���ˀ?�F�H�Ob�E� �cXx��Y-k����D7-?Q)K搹�%�&B����<����&���#c}!q=f������ٍ@^L��+��*y��'�m� ".f0�K@\�x�
×�3��HѶaCW��ȶ�8������ċtN�?,��a�����\|Rα�J\ʥ��rg�B�Ro�_�V�^��g�`�ۏtƶ��,�WL�� MtFaǕ��g=dls:�<�1�9k�A��`l�tg�*��ɲ��O�-·�/d~�A�E�n_��s��c�Nzm�������.�����s�(�@ɇ�J��Π�{�mP�,ļ���{�6I1(���M�Z:���K��<�b�c� �G�C�Iz����C���6Ϗ[�Pl*����.ǔ�s3��K�U����@�ό�$�)�!��~`*�Ω��|j���� ��n:S�M��6󒞗<Ny���� ��{z�o�/׃j]���g�6g�Q|�H�,$g?��g)�1<��ۑO*#Ջ�N�l��]:�e�h�,��\�JLW"���P\�2w��r�S]��"�پ/t2`.`U�7�'=��x��eO{��@ۄ���D�6/e`n7��<P?��O�Ȋ�����2�Dw��b2��?����������H>A�V�g�ɬ&blr�3��쓱�*[烁˰���)J	����`�'�	Lp-��=7�>����_6;_�����Wѝ��"��IXRƩ73s?5���N��{Џ�T���"e� YfaR����c�d6K�i���y��<���m������0[#�y��b:n���NV#Q'}�>mH{*�Vg= 3y��u��K�q$�w(Sm�T���^���!J��.7� {`FW���hS����{e��R;)dz�-��kn}}�`D�+�Ӊ���oQ�ə��/�-p���xn���c)������w�7��yU��̛dk{lZ$"~5��Jɫ�큜Y���w��I�J�h��{s�[Kۦ.�
�iW�n�j=�e"��8�&X
س�{�25���s�г�n��S2�����N���]��i�փ�?-*@:2hޟ4�p>�����/�=�C�#��Z����Ko"=�.�+�]�Z�`gڌCf��*ou�`��"����pz4q����i�|��ܝE+o�tcʉ�-=� L�&I��
�U|M!! =<`���C@� �7��I����O�Xk�����#0)�$�������x�e�W���0�Z��m�#A��h��uّG4n���o�y>R �0��U����!��/� 2�k��������1���%��F�X,��#���Y���^;���2#ir���+~�I<)�q�hl�F�4��r���t�B��v[�U��Y>��a�����l,\�g�����(��s4>�d�#�T�Pc�o3�ۘ��+9R����^J�D��F��eU� �����ܽ�'l*\K��G��s���ŉe���*�E�7�6��?�I��r�o��<�We6Vl)�R+�L�Ym��?���D���$e��xҾD����L,��
����������[,-�yT�^�@��zbj*�'�W���f���g��O����M� D4����x�]E ���6(ͪ.�`� ��J%%%٥�=��Z7@�;�w�ś���q��0ȷ���&�9�(QB�Z�ѿ}��l�H�%/��:���T��1�f�y���w8�:���IB�9����Y�&�F��%�Ŷ#�eog}!�n�|�A,	S����
[q�\��S����4� ���?��h��	k![������m�k��lG�d5pI�vYԧh��͍���^(hY���jC��k5s9�����؆�?6�[$z���ª�'jO�&�sg���==�LR�V����a����mhg�\�*�܄�������ͮ��P����v
�׿�=��7.T�ݻ5�U:S{��EĐ��v�P�[�و��ا�bd�b��q���æ�LH�	�'`#�o9�����;��������b�\�z�m*�������p�b�߄o���nC-<w����]֟*6Ə���<,c{��]��f祃��w��|C���kN��QJ��ww��r�V)��*�'N�/���iE~?�OOQ��d��	�#k;��+?��,-��E[��B���
=��8���C[�+�:�����}Ru<�K��F�a�8p
�]z�%�!��)��i�!bxs6��X��am�v��ַ'N��D�`�?�1���f;���bC<G,��T��Q�����Ym1�R�p�����_�z��N��XP�
�S~�֓].��F5���Q������;o�D�
<.��Eǔ�a�F��+�J�X��w_�AhAX͡�y��;����J��m`g�P�Q����v�@2���w�������&ϰm+�2��?n��>��]G_���*���d�_?U��#���h�Tߨ�u�!�GT��L��#�E�h�^��!u�����T����8���v�Ŝ*e�p��i��!���f+�1��0r؃��!%��C&���e<�u~���s��a���h�ܢ���u���UM�'������|�L�S,-�0���s[���?b�vC���Ո����D��U�@��09p�bx��Ǉ�tܑwѡ߼.�����r��9�	��@��8��)J�{R��o�a��sN���-{�}w�hω�����E�[,m�䂈c�od
Xp҆�u}Y(�ROGy�p��t�{cm��k��t�tq�@=ۼ'~%�'p��I��K|��a4 ���,u�W)#=f˳1�%�a��k��Ę�wM���'/@�ܡ��{C�I$� RE�{�We=m�i<;Ψ/w�_�P�@Li$pK��w���I��Y�~7���	=�^UT6@^�âL�Ba�(�ć�@��~s��c�獐�FA��W��y5�`��u�P��`+����@07�7�%�M��zrj���:��2π��楳a�j+�w���v�hSWU ��2�G�h�=Dת��%��E��E� s8�0?��X�@I�Y}�+䦌�ܮ1|ʂ^@��� `��W:G��Yd�n��?+����M��3>K14�c�����]���<���@?��	�[3_0��H�����D��H�9N��s@�e�[�0�m1�5���{H��qQlҕ��߫��ލ�7h������� �ʬ|��Kx���n�>�z����Y"C9�mx���
�(�E�M��5����_�|e���N��V�jX/���E������4ě'� ��QGN�]3�`Y���g�����IN[��0<� G��.q���u[s}��;4�\(�����:����g-ƀ��h��u�::p�rG��F�N�O&I<����F��g	���锳:�\�|}:4O�2:T�x�v�[��B)w���`\������НW�T,��)ݼC�`)�>�n�s���}zv����Cn�+b����&�c�eK^�����r9%����U#s�	��BJ��5��u���(�j�lK�f��;�����$�j��&�\�7,�8�jQ��ρ�|Gm��K�P妘w��$��6S	j�{Hn�u�R
���m!i){;V�q5c����\��$֩)�c@�9��kJ^�lz���D�0d�OP,�x��'��k#�6�)�m��|���E6\Ć�?Xx+����u�
�Oi�o�|v(���?EIy_
u�Fr�w���������m7j��N����,;��M�p��l$�Uq�5U���q�Rf�����,E�r������ǝ�5�P���C���^	>�-����J_��Ӄg�����k�'"�C-��yK�<Ր��ٳ�D�ZX��%�����W�˞$�#����e�r�.P����:�=jJͭ��r�D���*~� ������:�� ��Lr���!A����L��[��L݌�E٠&."�ha��X"�j|��359"�&�l����:oOl�^a]e��[	3/��{�;-��<�t-Ӹ6� /4�u��HT���J;�����j��Lc���V֡�H�S�m(i�/OT9�	T��a��J��K�91���~S�S-9��4plݢ!���(�G�S����i� ��:�(���I�vA�T���-�]�����Y�C%���*�����m.�RV7����ɴ$Q��H-7L�F>���c�V�Z1;9Uh�^���
߰ۆ�Q4�o���(���՗�tK}F���E�)|��b^�BQz��H:
׃Y�[�}F	BDe*O(4=N��YW�fa�j��
��o��N����yd�:����W���\0�\��`���G[1�l���Z�dk,'	���n������%]=
1�U}vl �����KS�"žN�)W+йb\�Y�^����I1�m��]{��MP�+(&�a4	
�=/�e�r��	.7qr*CnS[?��'K������~�Lq̿�0@�AQr���k�;�B�|#�d��X*��Tғ��9Ćrd��P��K�(̠Z����Cq_f�^�X�=;B�&ޯ+����O��E��k]��p��sɚgt�Pc&B����8'��Wt��:H!m2Rs*���{9;�V�h��N�M�GЎ���X�?�k�+<yfq$u���?𻋚 Mc?�#$'�nqx�'Ь!���_�ő?�'j�g>u��ߒ4x��UaKm'�.B,M`�yN�R��n6e>��h4
���S�#�*
a��#��Y���m4Et�F�Y�L��RM;��2�D�p�接��sZ�V�w��+���1�1qt�{.`�:�-����M��F�.��~���Dzuߩي�[B!�#,�q�ɗ�z�_���#�C���re�B�|��vT�]i��
�Z?���2��j���c�Q� �R�i�ס*+圁�A��n.�
E��D�W��"i�����39;��%���VC}	Dw{A�xa�ۚ� R�'��PYkZ�e3�C=���[�]��Tv��|�R^���PGT�u4:���	Aa_���q�<��e������t�	q~���"x�%��lU�`5���[�;ګ%�w/�'�I�)JIŵ.��B{Ѡù����i�x��鄖}A�u�Ef^���O���}%֣{�`"V?��UP���&^�,)CK!Gpq�cg��zY
0�n�^0G<-��뚼1n�!y
�4�a�����\J8p���K������tm\Jy�Wm��V~�e_�����h��wm��$xY>��\lvA�&km_GFd@���t��$�9��4��E�l�q���N�ݔ�n�k�'���9�X>~o����������o�P�k�c�<��=p� 8�����}�|*e$%@$���6��.��} ��bE�����X^�z[[��,�qN첲yn�d��bw����YH�%�z�N#�E���]u�+u� �U����q��j'���q��ЂX��R�ˇ�b"޺ԇBy��}f���Ee�.�+)�o�V�z"b��Ξsj�>���{8�6|*�.������@�P�_�@q��wo)��f{!l T���/L�����U��/�)�+�u�ѭ)�����y�2��N�H�0fUߨW�!E'́�&��/׬����[⮯�G�j��zp�w��<�z�]/,�/4)�4��恿j���E		�����<�66�k��Ai�����Rf�����	��@N��Oۉ�Z+�\�������N�&?K{��������Bx��֦u���2�(�h��5� ��w�F��_��˲N�d�PMY�$I�m�J�6�+�i���M�W鏣bю{�s�(!��'J�}G�F�/\x	�����d�W��9Z�m�̜#�b���(��uq��
2gEi�fi�I>�b6c��0���m�s_�q5�h��UwC9(§0�K�k!L'DW�)@k�l��e/m�>XN�����mK�HK� �����	\�	�%jf�	�Xļ�}R����"I!W���a���%
J;�Q��� ��
y��p�����Y�o�ĭ�tc�˂�k�-�:�;���Q����}>��\�1Tx~Q��B�p���R}�?"f�c@�@U�:�(�8��*�m��TFִ�m�f���KM��xR�,��>�5��aЈ��^8���Ę�^��]	�`x=�����RGSϱ��/�����_����PR�Fc_�D�^T�Pg~<�j�����,SC����t3솕��lg072l@zq���f�FҹAaA�l�t���̉�����0��f/q�oA�g����t�8Ғ��>I�q΀�ѳ��	����(�tB�c��<�2m���,�Z)�1�*6S��(�ߍM;7B� EO~���|;c�[���P|�����Ʌ��h�ϼ�]P9��|���Fєh.�3��;�B����Ϲ����2�!-��`7�©^��jHS���灛^�ngX�M�9k6`���I�é�`k�M��{g ������?��j��6���^˜H}]�g����T9�1����Q��%��إ�y��]灆��_��	n�ז'"*����qi��m��0]�jl"��/a|�.���7ΠҸw/�}=O�����"]�UwD�8e�2D7��<[�� �`ȗ]��65�0m�Dd����3G�H��ɵ�;�Q�����BKVP�����b�X��`���`����*���`��RB�v~��s(��A?��Rp�*�=������������Q���䉊����YUR3��3�v�ş������h�?�ᩮ�OZ &�R�M�p d�����5�����A�򿤳���O0hԦy��W:��P�;��Q��>��dH�o� <gJn�y��}���+Kv@nʥ#�S��T����>��.u�hA�7�B�`3�!��bS����H氥�Փdb�-���nʜ�`1��`�����qQ�$�6Q|���-��Ŋ���	��EyA�r�D̺�My�h��H��kȅe 5d5�]�y�YWצ����������-��[l��(�[l��6̞nByN�r�%��C&�2���;2��0�C@#����nn�3S?;����3���"�J�Ri�.��lve@�K�f�ƹ�����|���0g��L��ZF�w7H"�L%�>ו
��Z`�4g���f�*o��Z���"J�&��@�4y �Jq�|��	��9Jo?�t0�R���n YD�I���
 	�|:�r!�����v픦��m�/7�+I��Ԏ�PaE�Q�N3�#]�$��ց��̜�����0�"R��ٞ#n���5�OuF�4{e<�;�>���0��U���/3x!�m�EXk!Ti�gO��j�����^en�s7Xт@�T|��3��cӫ;=�����b���9m��)N�mhy}���R�r��a�����v.F�Uc��>	F����jV���T�eK����翌�A�>�#�ɮP&No�����rv9�(M�߻Ԕ�ݱUF�S��e9�1�c�� �u�*��+�S���[���e5�*�+37��^6��?��T�?��PaWr�|Wߣ�@L�m�!?"�|Dm��q*�	��I6�D�L�.�%2��?�ս���t��S�&<�^�����j�E��M���fo������v�}:ך^t 1X֡3�����x��E��_����W�$48� ϵ�%���R���
�oZ��6;�r����E�&;�7��f��(u!Z��{����l>�ir ��4jէ/����
�3pV���8
���yB��� PY�XF�e6%P�x�bmot"���Ǝ�~S�$ғ�[I�m\W�(\}g���O [h?%HIhsH	�0_[�p�`�����lT�5�v���h�E��^T���MYq�c��`���أ5 fJ�)��ŒF̿���<�l-��R2'�t��Z�s��z~�=$����j$�aص�z���	���)A�x�~�~�R��?v�n
�v{~�̪��{$.�H��"��:���"^��]�v/�~[!�S��O��J�Occq,*����HO���|��R��ވR�н|�z��b5��G`**{�L���=��b�oܴWn�$�w��*�*����$<�}�fJ��}�5���w>��|H#�{pR[TQ���!��_��)SZ��������g�?��.QV)2�#�o#��+��N!+lH!,ԲR�r����o]�e���qy8�}��F?+�S����}��c<�S�ƥF�g8]�r]���N�G)�C����TsC���i9�. _�c,�D� �\`Y<��>��so��N�cC��I��Y\m���'��&{Q1_Gp����T�(z�IE�����Q~�M]�xxF��]�����`���1,
�4%�%������F&/+��X���wd�.D�A�&��z�|,w�Z�"��mlk��J�l6� �2�FۑD������3�m��[2�w�?[��>)��G��w���|�	�B_L'�47[��7T�[u92�G���L�]��9��kD�!"�U�HYT~���K�k�&v��ig��"v�!Q��fxH��}2re��N���خI�����0�$߮8.�t˩ijB��.���bMf����Ւ����z<-p5Ě�	�j�bL�C�)��5�C�󖶧O�}踯m�0I8b��lǔZt���üc��u#��J	ᴣ��v�@��݉_�mJ3�*��m�ap�:N��P-He��4�w�"s�v��J�X[ �5�q{dc��d�i�����h(>�MGi�xp��k^��c9T��h88��kt~�(=�r~r �pۥ��L�I;�GaJ��h��dQ=ޟ~�����B������>!�0�t/M���N�x{��$��E"h���
��i����<��P^���0$]�q�@���f����~���e���6��NÏ��B����n�O~��]c�����t���|�Dv�y��*��P�M&�$��֒������:6���ZLjԝ�+�2<�i�V��`��jxK�w���vvѬ�& sS�2�8@�u�?D�H��r-��
7�>�-?��a�L�MM"|Y*��X4��t61	bb��t�Tσ�/��GCXY��?�+��ͪڏ�3k�\4�;��S)��ӰK���.��@,�Q�Ɋ3�s�B��(��D��ÞbNԾ@
��eU�V�]�1~[����{U~��.�� �ߘc���K�4�h�'���v�B�)aKK�Z-��ٮ�k��F\�&Bo9`�x�-I��E��!������}�І���e�#N+��w\���b"bg��B7wm�T���kKN7\�3$@h`k68�y��̓I���]�� �z�󞗬�Qu���p@�IźM�:$�d{�3C�u1�uK�~:�RG��[F/HQOStPП[g�F~gz??����\�6�}�j�O�:)T��H��S-ཤM)�b��<�\�T�bP�����!�����aPQ�)l�n����a�zr*��NQK2��,�����ӝ��,8K���o����IFU/���z�ݽ��\ek��5�l�@���*7jV��KP��}��&�WIɮ�Hh�d�G8ގ@j��}ώv2|�nG���8���3=���Z7�	�WCH'$�"1RW�m�ZtOi�\6V��50*Ar�<��ב�k���@ac-�O�? �kwNPlGzbN:��|0*�O�@:x�zX�'pkP���`����N�|��E��z�.Q�x�W�*N
���i�	��_B���E�q�
��_��L��;��a��9
\7w��乣Q�\��,(PM�X3\�$�?q:Y��T'�����,2ɑ�zLþ0�Ɇ����PM&��n>i����O{J�![Ӱ��ԭ�N��%Mk�2꘾����{B�)!h�H�t�q�4X�N�%�J-� ~L�xh��p���-�k�r��ѷ��:��8w�[�s5r�@ ք�~�4�כ��s�:%`�����L"��n:������\�7��^��3��\/�qaM��"�`��y�9��/&����.�x(�Oy�Ha����KOR3_b�$;Z}<�F)�$�}�ů' ����~�HA}�L�Q;C��m N��4�L��~�V#��H���m��q�\Uk9^�K�`���W�9ar�چ
署�����8��p9e����P״�S���Va���U�u�KAQԭ��2��
�z�F���0�;�SV��#G7m���V�%,�7��a���u��S���ۣs�%��#�V8�;F�Ohi'���/��.Q�dq�t�(�Q��|�����K}���E!������@	BF���t^
Dw�       Ĵ���	����Zv)C�'l���3ቍ+F�h��aj@�O��dU�[6��+B��iwV�[��
lrYmڑ�Ms��i����%���!V`S��T�>:ӏT�M�:�v�:<��#<�Gd���{�G��/S$��eѾ ����
�<�FE�Ev7퇱��9O� J�D��fT� �jd8��
�6��{CP$D���
�E�>�O<���&����jN�w�>��ի�qa�y�0�IO��x�6O8��G,NiOf(Q�#Ҧc�6���|R,Y�'u��%�D @K^���ip�
�u
lEBki�����i9(��dIO�����+gz mF	�*���^�O��3�O&�*�G�ތz�AM!y;^]���>���<�H\�➬�R!�9fg�Xk�蛩V���b��eȈ�:�O���`��)�8��w�� B��Iq�3�Ob�J��U�������񃑭!n�|SRΟ�����O�����5e�|A��0~���i���=;`�Dx��s�'��	0h�.:Iƾj�|e"�����	�O���N<y�s����W \=FHR&Qd?A,7�~�<�r��M��LJ1G�s�R�F�ܟ��O�����fӖb>Ź¥sݭ�;`��M�ӈ�yG�$\�c�
u�=qN+��>�'~]��ED0����/Y���1��>�A�1n>v"<IC"�|�`����Yd� �CNK�<�Da 2  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                