MPQ    ��    h�  h                                                                                 �M=��ʻ���1�M�0���K<4u�۠���E��?w�����`�l��<�+�����R�W5 zB��ִTk}X�I�e��A��R������[B[��r9\eX1�j�SHgT�[�3���b'��0�~�Fčޔ�;�^��!��iP$7E�|�E
�����W�6w�~
Hc?ܓt54�`��d�R��oT�4rǒ`d?�Jf��8�ߋZ��$�G
��&�}����a��	IgU%s%���� Ra~+7�@vf���K2a���~v_8������Ŏ �����'�N�l���j�%?�j6^�t�����I���u���WB�x��z�p+-Аn���7��V�r	�.��#�k��N�:�'�佐�f4T�����{,D���B�JZ�>ٜ*�z�e1�k4�����:x9mPn�Rq�i�Rz� ƻ�ێ.����,��hwq�`muW�<&�Fd������Z>p�.q_�ڍj0��q�2(��t��gޑ�C��F��
P#�(2��*1!��=P7y{����g3�\��`����q�/����!�c<��k�����I� eL�W����+[
��L�!�?_`Nd�j��((�� _�U�ً� "�Q4�W`�4-��p]v��E8�|�b0��_�<c�qvvl8����!�9d=����4��gi���&$|�~�4'��B͞� $&ؓ�$�ȝ>��_�)Z|�8f����jNB;�FO?��@������_�R���5DqY(�S3����(P�4�������X��Qe�x��˳�h��d�Í��~���
e����
OO���&�ZV�^�[�;ܷ,�Z�����t[�����Ċъc����| zoͩ���/!R�Pk�gu��"+@�;ψ������=y�ٽ���?�1f����G����}3!��dߚ^��ۜ���qv]E�i�Ż8~T�X*R�#�j���[W���{#��Y��,$`bGbh�\�������8�>�
��Q��k8�Nxg�Jy6���t�R�K�
N��P-L�}��,�R�*�]B!jg�Z�w[�nS�1:��we`F�8�8�:X�{�FoЉA{՘9�i1�mY�p�2��r�O?�9;�SL6bW��~&��Y?j�uG�1��Q7���\��XO~D+�b�z��8h�>0NPލ�9�a���pBvP�)���@HWV˻'*<�g��>$�ޤ|{�n@W16WMa��	�G�����^oX4��'����jR.D��u��x��O\��4�9��HS��U��^�xf �:���k־�y���`Tn�N���	5��%�5�����L�	8u�����'�ba*�������ĺ�W�u7�Cs l|����r6b��bx�k��y��e��3-��?�,����~���;�����0�;o3�F+�����
���N�E�F_��PL��`�Z���g��MB���ʾ��(}v���b���;Cv���[�.n������X����J.�վ�d`{�b��zwM8� �����2|��J�? �pׁ1rh�%U����е�CN	�D�׷��^gK9(w˅&FH܄������^�,z�a˔��Z%<���:Ζ�R:��>����m�c&P��]�p��lH\+?J�B��o�;�������a&U�$�����07��'&BOC~t�$\�yJ�a�6R]�i�o��CH��5��w*��ld��_ٴ�;"s�0�$HۑJ �&�"ǯ5Ւ��q
΀�s���{�m/.X��m���'ñp���k4g�s���-��cA���]�m���+s�uWb؟�D�FU7�!�&}.b�*� 5,��}R��G��O�I�j�X`�^��nD0��{��%��J��q�E5d���s����5�p��C���UDRڲ(�����LF�1:6����'��tP�.�؅��!s�0��N�h��F#�~Fw�{�hY�ک}����*Y�<,�ľm�������Μ����=+�����D���Y�E���w�� ݨ����nY�]+�����<�׸�Ԃ]
7H���S�M��r.w~�B�c�Ӗ1ư�K����aht�Yr-/��nX�K�߿�<��a���[���r��l)��5nbv�Q�9�RFY^H�������)�+�l%�.�V*�����en�����
���LB��J%]�bs[s��uX��1<s�����Ѐ�OZX!��Z7-� ���Zĸ��46��V��i��@�]7_�@.�`Gl&��>A�F��y�5�-��$��C"%&F:nDE|�}go�D,K� ���Xn��0��2^�k�c�������H4��h}�{���7j�RxԗD��J��V[Q85�m_������,"Fq�DTM�VG��#���rP��0�����
��W�f� Y[0h�E�Ӣ�~�V�@_�|�.�"���*� �t�r��/)��E���Ԉ��<���{j0,�e� %y� �J��A�o̡�%U����1p@|��g�VXI�ӋS��ڔ��?�5�FL�H^�|�����"n���T��!uc�("��d��"�߸�#�^�Dbi��Vm42�	ߛ�� %��R.���:f}c�6���)ݎ�gg�S�$rl٦p���l}j�$N�����t8M���.ܖa|�Y�ݫ�k����z���a�!:ْ*zE�t��,��Dn��g:G��4ڿ;�)��y��fs��y��Rh~l���*m�v�	\$Z��-r�]&��k��.��$��[��o�h�j��"3ɹ���Ƞ�FS3��`���6�(�~oQ��>F��|����;��Vpi/�b����4�қ2�ӟJ��Ԍ�1��m[`K�2�1h!r�@��B����d�`�۠9�<�X���x@��6�G1��!�rT�VU�,�:.|�a�u�}2V�I%�
zV"*`d(E�W�93�yo��C@��D�=����/��iF-x��U��e���wBPRÃ�Cð�/�,���%x��(X9xC2U��q�푑�C{M�d=7<���/mV�0G�Z�5���@����<v��FA4B�P��{Άmwfx�(l$�غ��9��b�al\&R�ޫB^��-�f���(��o�ҧ�\���/��Kk2�ȹ�f�|��I����}]�r*��(4B��R4T>L ��1s5�@� �H���CܮM4/�'�ϣ��&a�}�O���R��#��N��&Ȼ�
���83֠��֢�/U ���'� 툆~&R���Eط�}K��� �v܎���@0̎����Tl�	�ld�j3���Eį�(�����Yf�ܖ�sx:z4'�-���-Fح��V_����b)#�*{N߶��b>��Xdf/�
�
3��m�D�(�B��,Z��e"� p:k/���Wx���P(�R�r�^�š;(x�v8b.��2�P�ˈ#��{l�W�&�
-d�X�y�>ka�q���%�v��1���2ةt#�^gyC�c}���P�.u(MdU*��{���yQ�5�G��ҥ�����`e����1�/0����"�<6.
��N���MIy��e�i�r�~�j:�
n�L��?� �_cj	��(Є� zxxt3�۪�Qo)�` `����v&b�8�R�}�JP���}�%�l�49��z�!@��=an��OC���X���λ$�V��6o�*MB(s� ʃOخVz�C�>����)�A�8}��ȩN�::>�
���w"�:�G�)��D1>�N�}��d�4�ˢb�Ѻ[8>���~��1ˮOfON���H�떛� �ey,a��}���h�&���Z�<[�>���5��e�9įM�}��������|!�ez�~��޵��jǬ��bl��}%���N�0�d���x=Tb��������fч��������3<|i��&�^�z�=*E���$v�7��4
�v�GT+Rz�ji��Px\�M��{�ʴ$ш�f`}��b���7H�6C���>�5�1�'�&����gs#6��vtӅ��晧Nz����y�8S�,�*�B�L�>��w��]S��	��O,`�?8ғy:ӹ%�!���|���\��;��\�p�����x?g���Lq�Q�?��&�Q�Y��wu�a���f!���\4O�Č+�|z:�8#.>/L>�}��@�a�eEp�'��$�E�g:Hf��B1w�|T�`�$Tv|�0{�i�Z1��M��E�$��Y��9T�42�'`vj�e�R��M�o�^�����9 �ZH���P�^~� ��z��f��jQ���c���cT	)���;	���%�q~�9�1�	c���X8��� V[�]=�*��I�~�� c���n�uRp~�q ����\�6�F��ʕk�$�n��iE�z6|,z_=�y�b�R����x�V�v���ܢ����E�����A��?-������u�4���LMQ����'��v��t�)Я��C��+���nq�D�8�h�k���?��`�y��d{�"b�kzR5��[�J���p�-�ڥhp��(p�&r��t%0��Q�4�Pp�N&i�2@ȨI�IfD]wF��F܅�����s�^�`���~��ky�<���:IP%R�	�y������c!O��<,pDj=Hw%JG@�J3�ǿۨ��8&P�ھ��h��k��B�O�]�O_\̴̓�f�6M�?i�D�es�x�@Q*���l��_t��;�ي�?�H�ܪ �@"B���mFqE7{��(����5�ȹ-X��^�'z'>����2�4�7���� ��AK�]g�\���������ND͌�7]/�!>�b
* ����o��q����I˻�X�=A����n�"�0G"@�t��?�L[�p|d&�D��Y1)h5qrd�^���РZڍ�R�N��,(�:�6Y�Q�	�5�zҩJG�˨!Y�0D�Ӯcm�F~s��{	x��U�m��/�e�U<��J�hA$�gw�������}��A��p���@̍�F]�@)� ZiлI���!����](���K�������eD���|�SR���~jH�S�p���,�)ɦ�:圥�t b�r�M�[\�̆�$�G��\����-p������1l�5I��ь����[^CkU�S-=���\+������V=��I��� wn�;ҡ��d�L]pJ�\�bNJ���?�PC@s��?�U�����X<xZ�����8�20G�N?6����JƘ�^;+�g_5�T.���lG���(�F���y<�?��\5$��"�:I4K|*i+oa�mK������X)Ы0�.`2ٹ��������"���cC�a�I��h8<_�,�7�t�S DM���si��Q��m&.�.�����_L��T���Gz��#��r�x�0�9x�ɹ
9�l�A]�Y�(�h(D���t�~Ph�@f�I���V��3#[?tc������)�V�ETX.ԣk�ҷ�5�V\!,����m�P$Jb\�E����v������p�1T��@��p�b�V_��y��n�y�\����,�p+GL4�f�w�Y�t��� Z�ϖ$�i��\ä��7�_SP"!�?��w¸_�K�%?m��	�	"�-��pk.v����
c��<�$CŎ��R̎l2$X��k�ǻ4��WÄ�\�����V��Т���ѫ����S߸�|S�<f����#E�t���𪌇n���ۖ����;�@@��}?fNE���&��J4~gT7�>���1U�\2Z6r�R�OS*�-�I���yҶ���*:�h!�j���ұ��U��;3FN�޻K��O&W�o�[g>!�7|�M���c�Vk�G������4Ǖ�2G��JҜ����nF^[[7��+�h�H�@��B�+����������,<Q���x�~��QgTG�t���Tج�:.w?WaD7}�B�d��
�>"Idc�W�<3�ƴ�l�2@�@�s �b�
&�i�
sxuc���}o�!��PEÞ	��`v��{',V����g��V9Ӆ�UWct����c*�?5�<��Q/�W+�DZS��X�f��=x�����Ao@xPWe΁�f`('Ȭ������l�ɰ��u�\���ަ�{jd�-�張�l�9�҂�n�Ͼa�m�Z2B���!K/�	S�W�-}8��e�e(�H�M8>�1t ItsPd��{/��I���,I4�#���HG�kC穀j�̒V�����<�������
9{���H������Uۜ��b[% �е~!����e�r��K�Lx�{yv��~�?a��⪎����1s�Ċ�l'��j�.� ,��;'�*�㓞*S�7�����x&�z��D-����hp��H��V����L�ϰ��?#"'�.NN��������WSf*8�^P�N�D�qcB[[Z{�������$k*ŵ�>sSx��KPC��Rg*G9��v�(�#.��ƫE�ަ����W�!�&�\#d��g>f)�q_��d��	�v��2���t^
g�"C��o�M�SP�lX(hY�*'2%���y�����ۀ�&�� ` e��7/�w��u<q��=�����I��8ez�N�K��ha
I��L$t^?�ZW9jdKI(�c� �.�ﬢ��S�Q��n`��1����v� E8j�^��R��l�������ln�J��"!��7=c$�jϕ�]h���@$�0�X/��~B�g& �}���Wھ2ˍ��)�&�8�	����N�Y\�Da�%�^��2�Tm�d��D�(�I�
�i=ƫפO-��݂��68������L_˩@��%؆�g�Ϟ��[�eT���d�����A&w{���b[�a��"�͆@Ij��=���<��@ڳ�wE&|<��zePݒ���ԥ9r�Gw��]�T���ɰ����K� �v��=/� �3��u��f�i������wHP3W`.�Z��^sb�x\��0E�v	����N�1�T1׳R�h�jD�����u��o{�&��݈��`�W�b^���&�qP��ng�>� ֌v����_�x3g���6�7�t�́TNu� ������,.SR*�d&B�O-�y�Pw��DS��բNHs`��e8�`:N�����#��-��o�z�Fb�#��pS0�C�?��	�`*L�* ���?&���Y��!u��U3	�-ۂr�\o��OB+-+���z���8��!J��F=�����a�px�����±3H͕#�]Xk2���;vc$R�[|;m�d��1��'M���?�5��dq�Y�4m']'��} �R���C�[��E}���.�9[/H�#�K@^i�� O���O��U�������3T�����&�	��%i�d�T�㲄��ʿ#�sG���>��X9�*;m2�9�	�!|�M�yu����$ ���#d6�"��;�k߿�����ĆԵ�,E�t�b��#��JŤ�qw"�<��r��䀌ׄ%J�<���)*�s���pT�].\M�������1Dv�T�&�j��C�Bz�Q��nL.֬s�%�k��� �a�46�d�[b�cEz-=,���-�Uj��(�8� �8��Q�p�ru��%������EN����������o�w���F�㴄9��'v^����R �&�!<��=:�)�R𻿔��0�.�"cnn�o:!p�3�H�SJ�k.�%�Й���g&K��Tʷ���*�]�WO9�J*}�\�B����6H�-i6��� ��O����*���l�)__n;S>���HQG/ �R"���H��q��\�U����6��#dmXP���B'�'�27���4ݒތ(H����A] b]"O��4<,�kn=��%D�Q7�\ebe� �#����Z���2�s�fI-1X��;��T@n�M�0���/��@K(�'���wd�ݯ�A%��5,���y"�K��h �>���	�'js:���a�P��$"��_9!�w\0�rЮ^zhF����o{$�=�Ю馲��s <bAi�c��NC>J��ƚ�3��K��{tS����;�o{\N�v�����P�d��]�ߌ�)�0���>,�q��}U6S!֯h��~E�R���1��'��&W�W	3t=yr#�*�6j���\����}�W�4�����^񀢕W����5$���[��ݕ^>:����|�G��+&����sV�ϔ�hM��4n��H�H�8�yiCLx��J|�b)Y}�*���t�s{5B°�m�bO�XW��Z��Eotةm%޸�ۇ6�Υ��V`3"@_��;.�
�l�]�t08F��y�L����$�_"�:$D�|etCo�	�K�l_�W
2X� �0w�2T@�����ÐR�'>6���Wh����G�z7`�.��D�1��5����Q��6m�l�I��"ť'ØT��*GUZ#��r0n��
��ͽ^Y�_h�b	��f�~���@�z3�d�w�j������ft�q��y)M�pE@~ԾJ+�2N�1n",)��6����OJ��/ ��@��S�-�1� �@<
�].�V�S��v[��W���k��������LϽG�r#����Q��;���J:��D�D�1Z�^mu�Z<"|�F�����zX6��{mꍲ	Un��AN��$�.���<c����|َ^����:$�cӦf���"����������j!�_�N�`�Ϗj�����B�#�;1)�W����9E]�C�"A��EnBn�����Ȫ9;�wx�o�~f)�6��?�����~b4%��ɠ���\M&�Z���r�gִ���}���Y����叧h<��j�Y�ؒ��4��8�FI���BF��0�(OcoGW�>�H4|G�q�cVf�[�A��F��4�x�2�@xJ������	?�[VCu��h�?�@)��B���Zg���uA�o9U���Êx� V�l �G'QF�~�TS/�b	J.r�a�v}�O0M
���"�!"d�	�WRF�3�3v�ǳ!@Q��<W�k����i��x����ߎ|�P�A�ù������,��w�[w��9.��U��#<�9l��M{<4�^/�+&��Z�0A����I�2���x�iA�^�P�<G�|�f��(�՛\��U�Ƥeמ�\\� ޡ��G'-�c���غ�"~�]�|����e㙉2�ţ��$�����	�}M���(jo�Hx>k� w�sk`����������$w94e����s�cϩ��ڔ����c��7%�w�E�\�ջ�
�
�Ȯߠ,x��z)�U�a�񝻠 #8�~��QE��-��K�	���f�v�N��z�mv�a���
)�ClB��j)ȇ��&��%��������<⒗���5�xA@"z*��-a�7ɣ���.�V�����"�_��#=�!�oMN�x���6y�k�f%�������	��D�0B���ZV2͜�(�6Mgk%H��0xjC�P^
=R�XG-��LͰ��[.�c�����X���KWD�&��)d>N�o�>ayqpFp��7p�3\�Yl2��1t���g�p�C������PT�(�n�*����G�y�dm�}�ȁi�m�`�M��.�/&{����|<�����YS�@8I/^e5G���6��`��
$�L_M�?0�Ukwj��I(Fb �6jFp��NQ��`V޻��vܾd8%Fv��F����^("�l	´���!��q=�w�̅{��ؗh��$-+���g���QB�{u @����d��9��\].),�87����(�NS��wo��@g��mr����쟒�DB@��D�S�ą��a��j�`�X���X����I�dˤ��Y��A%�!'���He/�49� {�����&�;+��a[դm��b��*�%N�lО��Wћ�!�2�Q|W+jz�A9��כ��u���:t�X���3/�K���f�$���:=
�o�nW��f�kF�X>N�2��3rd[���^Nن������ޛvd��z����TL��Rp;�j	�����t�{( �j3
�]L�`�1^b���5�����	׻>�c���8��h>=g$�6��EtIL��/iNp��a����d�,Iq*B�r���t@w,$Sؼ���`:`w!8�N:ɖ���x%��˘
�'�
��~Àp����C?]%���L�b�u��&�OYPU�ux"Nz��o0M�x\�3
Oݱ%+��z�-8���e�V���ʽ%a@��p�L��s�v-H��U�x�������$��U|��C�_�61G��MJ��Z�(�O����}`4���'���x�oR?3L�F\��x��=����d9���H$V`�F��^��� 
�>�5W��a�i�\�:�wT?D���wd	F}�%$Iϴov�����ʚI��(�VG�SUk*����ƥ�6���ȑ2u��Y�o� =wޞz
76s�R���"k��Q�d�y��@���*,����o>��L[�ⴌ�+6��H��M�h从��o �7v�E��.�K����ذ�M����Y��]�v�]�*n�%ߟC��p�̈�n'�����)�(����[%����wd�z[bw|Tze�ѱd���ϋ#���[�a�p�p(B�r�2k%晦���pІ;uN�W��谫��y����w<1�F�ay�t?/ܩ�Q^�(��rEV��<���:?#R��%��)\��p�c�{��X�p�+H�.�J�h� �S�=>¨��&F�Z���a5C�x�~O�\S��\B(��2��6C|�i�\����GVը*���l�1_�z8;�>�A^H�� :m"8��#�`q��q�������ޖ~.�X��]�v'4�L��4��*��.�A�H]��A�O�d��)�i�lDCy~7��" ob�+8 fO��Ε��g�׭Nq�IA�1X1�N�� �nU�(0�o��Jp8���=�=���'d\S��,���5��2Ĕ�r�ƹO�CL�y�$����"̳:GY��-��k@ҟ�h��6]!�)�0zlE�Y�|F4�KwC{?�{�K����0�<���^��F%�,Ŝ��O��Բ&���<M�|���6���~s�1m�H��R�]����d��'���]�Q�8NS<B��}~ .�ɝ�����"q�\����^t68r��E��=��Ej�}��R��l4���mր�{ނ'�'5����P��#Y^9)��	�|���+A�Ӈ��:V�$u��g��V�Jn����b�4��L�]#J��b�j�J45��ưsv�������Xr<CZwv$JN���:�����6�T�� EW�Ԑ�N��_+a�.^�l�&��X�F�_y���^Ȥ$��""�':�sG|���o��xK�R�����X�Q�0/�62�p�圓�V*ِ�}�9�ܦ�'�h�Ӳ�bR�7��#	�D�r+��$��j�QI��m�ӄ�dN����JT�#G�(\#�a�ra��0)�����
/&{����Y�Jh^����x�~�@����X�en޻  ��t�����V�)�/5E�G���I ҭ0���3,dM!� ��J������*5�.T�Z
�1�x�@ך[�X�XV&�z���,��R�)�vwK��DLj� �ma��P�Z�Vg�����ҿ������UE�"����T���)�"�m�k�	��X�����.,qJ�kBcј/���9�9���$C�$�a#0�}�	�U�3��>����c�:��Gl�*ë�I���H���r~�~��E8��]�p��oun��Kd��e�P;�8���If9i�*�#�~]4����jͧ
�\hhZ!�r]�����C�cU���$��l�~���hW]j�)y�rs�3���q{�FD���q���g1NCg�o�r>�Ӡ|X�D��Va,l�s�ƥ�4�{=2=�vJ�腌K���W&[Qo�Cb�hRV�@Dz6B�n�5HB�r��
���	����xq�����G�M �
�T�Z����.m�a��}c|���
u�R"�X�d��Wퟨ3����"�@��9������ɮi�$x��H�����P��%������u�,�ӂ����1�9�j!U��E�>��ⴔH����<oϿ/>Ǝ!�^Z	��J��5��pܥS�?A�(PTB!�w8�f�t(�o��)l��yJ��q�0\�C�ޜn
 K--?�ͼ�"m��+��8;X�b���82��8���:K?�M^�}�0��q (��C">]�� ���s�|�q0@�rG+�_�4 g����SN������LN֪�q��M�������
���i���Gj��^�U�FP��;P ��<~c^�e����K�毧q�vm���WK����U�e?�:�l]\8j��͂�a��`H��`]^��,!���+�Cq.x\�6z�
�-<hE�ޒ��~� V��K�WY#XCYy�xNp	x���)��f 0G�=��AD"dFB��Z1ni�����k �6����x% Py~�R]���-I��f�G�.�I5�a��TV���)NW��
&{`@dyּJ��>\�q�M�V*#�}ml�2�.�tԬ�gJP�C�|���PH�(���*��ݩ/JyH��QU����q�`�VO�I2/�����{e<瘞�s����I��qe�ڥ��AF��%�
�:�L�F8?�"P��j��(�� �����i�lQ �V`�޶�tv7�D8��Q���d���֨�5]�}l��v��x�!Q��=���̠G��S�c�q+$hE�T���B9�� �b����ڴG��7Gf)FQ&8҂ն��N��:2��[	`��WX��]H����D�w��?Y�R<7���'ע��E��8�=A���qB˟ч`g���Ұ<�]��2�e
��tQ���^��K�&-�M:[�Y�)q��T{�`�o坞�4����/��!|ry(z[S��o&��b�}��S��DT��f��q�lX=�n�٩ns�L�f������A�3����P��^)p��� -�f�v�P���y�ŧ׽Tg�]R�-�j�D"����K{����V��`�+�bTQ�Ȅt��@���fi>���BW�W/�2#g���6dG%t��W̷)�Nk́��C�i�,d�w*���B������w�y�S��a���`2e>8#eE:D�k�f��-`���n�����&�pɭ���o�?؎��r�L"sy�1�&���Y��u3|�i�#$*(�\��BOxXv+��8zK�.8T|��`<�ť�]a{d
p��;�>E�xZ'HCU����(�c���$�sc|qF�Z�1�ԻM�-�u���o����4�Ǫ'1��s��R�m~̸���;���9��JH����Al�^NS Ž6�P���J�D%��uy/T�Y����	�%%�佴��_�zf��u�a�)��o��N�l*�������Q���CSu���/|� �
[�uF6ΙB�Nkr����Y���y�+?,K�\�jv�&��������2�{�( *����׺�.�2P���w����+�SSM���锿����kv��l��?��1�C�v�Gv�nH����;���������ժѤd�$b�/z�`��﯋�Ë�.ڶ@�+�pC�vrk��%����H=�!Q�N� ��C�ݨzm
�%-w���Fm�̈́���DE^��_��X,����<�Qf:�<�R�-<�*�;�d\�cŲ%�Kpu'HH�o�J���ۮ��x�s�Re�&A�$�
}���?�O/����\}���K�6>q}i� ��.^q��&*q;lP_E��;�ۊ�7H�|� Uon"�����Kq��������,͖��X����x��'�3.�Z��4S���^-	ꄨA+�]��J�j̅�a�D$D~7.�A�bl� !�v��X���!��)g�I|o�X�gy��0n�l0xFf�e�6���E1E�d�D.杏pB�W5�7@į4,�Av<���G2GP�NP:�?���І�i��\-q!
��0�2�T�F���2�{ZeB��3��h�1��<�*n�Y)��x]'�/
��.5�)�d�Y6��${�̴�1rE1����z�+J�Z;j]������Sf����zkv,��f4SWN��^<W~��#��'AvU��}ɷ6��0tQS�rim���T�7Ok�?��ME������^�_�؁���h�5څy�=d����^48��d�<��PI+\qH���MV��������n�iJ���l����L�9J�b��G��^��!8sq_��fV��� X�uZ� �%HH��oH�u;6��3�[�搏�6if�_�V.94�l�f�Ī��F�@�yMaߕ��$z�"h6:��=|��oo2OBK�X��u�XZ��0Jg~2J���w�9���b����4��Z�hi�"�}�Q7V��䫙D��X�k����Q��RmKZ���V���D�T9��GK�#��Pr��N0��E�
��t����YG.Qh��[濪e~a\U@K�z��&��ޖǆf�t4�P�|S�)��E�o*��h]�(3����T,��ll7��H{JsR�vL}��4a�|�51�@r:e�S4�Vp�5��!C��|��QS�!�@L���h�Aj�Nǅ�qG��@�d��b;n!��8$�Pn�"2A�����#��Pm�i�	�����ז��].��U�&!�c�N忕O��K5�?Yh$�ڭ�\����6�5���߽�`��0�܂��ŷ���ӭ��OM�������ڒ���E���� �{� n�l��X�� �;!F��e-�f�⫤e����)~XTձO�T�b�\���Z�Ɠr8�F� Ğ��LL�����T�[�`hr`�jy��rL�n�����F?K���]�"Rx^�Wo=�B>�~}|� �ԧl�V\�x��ac����4��2�-�Jc>ጆ��?��[L�w��-Th�c@_�B@z�I��L�w��`N� ����bx,d/���Gj���T�3Y���.h�taU;�}���
�W"���dN�W�3�mm�}, @�g�T����͛��i2b#xF�t�����2�_P>��������o"�,��?|t�9��U���Yf��/݉����<�"u/ـ���Zd�R��1�P���(��.��A �.P�g��r�fq�f(Xs��D�������ZZMQc\��ޗ|{n�-�`8��)�wU��^�H�N2^��G�2SB��R8��U�!����}�4~�;(���>\>�=� z��s������j�M��ܚk�4�8����>���tI���Q��X�^˟���ߒID���
J�=�$^x�b|��p�UlK���3 Yg�~��EأbK�w��kvH����}��W�����A����TlxD�j����)ě�ڷ����]�H3���xw�Sz AF-n��TH��7V�]Ʃ��=\#s��R�NK���N�@���f�(�o��t�D=�B`�Z�՜Q��l��k��O��x�DP�R���4U�'���6.Ҧ�Ƽ�2�����W��&Vgd�Ӽ�xn>WA�q&ut�=�
�&甍2o�zt�Eg�O�C�o��^n�P��(��1*���݄7y=K������݄�#�Z`Q2�drW/�<�h.�<"�����2I�Ne����l��V�E
ژ6L�_�?fc�K�Gjue+(��! ��`ُ�G`Q[�X`�N]ޱːv���8������<ֳփ��"l?ϐ��b$!�ȅ=M6̻3���V��L�p$���|@��=GB� �B�� �/��Q�)��o8moG���N	x��$��v���c]m����JDx���:j�z�<�,ˤ���NZ�����x�/�4�˚����ط�W7�ιe�����V���,o&���FY�[�L��Ն�
\ěg�}����l�Q����|��zքu�Jy`�VN��"�N����9������u���-=�z����c�F��f��H�!����3���˄�^'T�)�b�r�v�]۩0&�b�T�Rf@�jզK�<-:���T{
��� �Èӱ�`�E�bϮ����"�L�?�>щ;֝�}DM(�gU�6?�Tt��~�RD�Nfzm���$�",�f*���Bh�*�{wb��S�"�_�H`���8>@D:��E�tىh)��@_���~�4��p����5�?S��+L]GD���&��rY��u�������of�\ �OO+�$�z��#8�%���;�ŀ��a�N4pI.������^!H��ƻ��x�f���C�$i�|�l�U��1��M��mܐ��E%��'4ȟ'��mn�R���9rY����~�{�9��HZ��<2>^z�> �k�����u�����[Tu���y}	��%��0���)�����P��$K�����I�*L���j4��lK¾4(u~�j�u s��p8�6)���	Q�k0{��Z��z�+�fS(,�m�e��X��{{���󕊭ޢg��1���Ubճ-�x��w��_������M��
��]����v�M��\�Л��C�@V�n���$L�_*y��!�j��e�d�Ĵbm�z��GXϯ&j���s�Ә��p^br�Y%��2�=�}м�N�	�枡��5��Ұ�w2��FH������ߨP^�pߑ(���W4�<�6:5v�R���eχ�g�c�J����p0Q)H�ЍJ�����ə�<����&<K�e��~ �bO�ۨ�Y�\�<^�h-`69��iGV��QBGI��0*L��l��_��>;	�����H�G� p�x".k���fq189�&GE���w�4#�X�5�˓�'*���5r=4�du��O\��_An`4]S���Ď�� �vKD��37ɥ��1bv�F ���<%�]hF�}�I�@�Xg`����n�O03=���������θ�el!�d��A�f��B�5]����-¼Ru��Z�.�o��H:��K�='UСh4ҕ(;�7Du!E�0����OaF���-�{u���A���Cw`�Q�<3�T�Tah�ӔIoRs���w����
�,-���W�,uJ�#~Ч@̨F����C�]r�{�����K��HUѹ8ட�Sr�үُ~֓��?���["�������Atl�er����S��rx ����H�m�"��대�d�Rs5����x���Y��^/g������x*�+w��y��Vq�0�5����~n�cաY�V��7+L�5wJ���b�E���7���sl$2���[���\X��.Zm� b����qy6�T1ζC��Jf��8�_!l�.��l3���E�F���y��Գ$$.7�"��0:�3�|V�o�!�K�~_�hZ4XSI0e�2ŧ��R����_�#�C/�H��(�h$�ۘX�7ю��qBD9U�V���Q�Qml��*���)����Tt0G�/#�OrR�0�@�*��
%����Y��+h�~���B~���@Q���zS����q��Gt�jt�wp{)^��E@����BңU!��c�,ڇ��2�0{J�9�1��^5��Z�$�1@�(@�&�N�V�*��/&��6��H5߶,��\x�L����c=����nB��Gu�������H<3�/�o�K�`"��\�ʆ{�˹&���wm{�@	�H��@�� �.�w���c%ÿ�����z=�$yFo�W���3���˾���1��n��ܽͅ�`���}��S92�l��V��t�E��S������Cn��Gm~�۸�;<�Q�ৄf������]�Y=V~S����'_�@;\�L�Z�rfǴ;�-��d���a�"�i�Q#h���j�*;i�u��ȧ`�F:!��'�x�ݒy��o�	d>�I�|�&��BZ|VWN��)"��w�{43��23ԗJ>�̌�����N[G'#��mh��@z�B|1���i���� �@$�W��V�rx�EB�`G��Xh�RT{,�35�.c�6a�|�}�5c���
k�"q&NdO��W#��3�:��ؘ�@�_lo�2��v�im��x�8��َ�,7P�i��
�8�F�J��,B�5�,f wצ9?�VUC�'�t+�E���T�<�~/t[&��Z���D\��k>.�o�	�;A[y�P����m
�f̱�(�h�_�P�o�W�5(;��)\-��ޒ�	ֱ-�G�!��Y�����`<�y���C2����r��pL�CgG}�X	Q�+(;���9�`>ױ 5efs��g��(� ���46*`����t��/n���<9�B��9Eu�(���-�_��K
�x���8{�}���),UGp��N�K �.�~��b4e�^l�K!�gH�v#^ʹ+�G햎�A����ݰ��l�LJj����7	��ԩ��x�����⣈���H�x��xz��	-��T5;ش�V���aݰ�D#��@o�SN&�����2�_f�f�F�ʩ��:�DX�IB�LZ�E���ԏ�?k�'��xx�9_P�ƀRSH�[Q�b�s�}h�.�#N��L�ʅe�H�WkK&1�d�伀-�>R�@q��&��o�%r�bb 2JgtJ��g�o�C�������P���(�m�*���__4yxn��NF���\�~�.`�y�҇/�Ey�C�<]���E��zI@W�efb������b�
�&L�b?ĊFg�j�X(w! G���"7�Q�>`'�ެ
�v�D8V�U�����^z��qzl���l�!`=vY��?m�I��'	�$��������B�xc qB\�5�ڪ�u��z)���8|Q���
Nd���V����ނ.�����P��DGu�5՗�Մg�BO����Ʉ:��w������˕@�(�r�ͰrＲ���e��:�=�����-!&�<���"[&.H�E�����֡�T6����!ѬG,�c`�|�uzQ�U�%�Jԑ�#ǳEv�I6�D߰|�J����bq�=�����(��I!f�1��i�c��3�0S�Fl�^����de���kSv��:���`�gvT�S(R�r�j�(��w꣟TB�{���{�P����`�^bJ,�~���]������>�L��?����hMg�l6��t�e���~`Na�r ����,��=*y�BC���e��w���S�gޢ�i�`�L'8Y;K::R,�h�������o����Mp?����?���]L�;äFe&ռYa`Lu���������y\[�0O� +��z��8ʥ���2{��[�a�XRp���(\�.�H����4��*�n$>~�|��e�P@�1XS�M{��ܫ������4Y��'g��i�RPB,�7>��?�1?��V.�9G�H��m�7�^�x� ;?S��/��uC��������Tݮ��*	W�^%U|'����p��+{8_���'!��Di�*���%�R��Y��96euY���� ���k6��b��B5kK����P��Ut�ԡ��,�Xծ`��]��6�=���(�����|�lU�����(�l[��_g\���#�I�Md
G�
z�.��v���;��V7IC+E�=��n����_�"�������l<L� ��d�b�Jz��ռ����T3���l��4)py"�raH%w� �xD2�W�_N��������t�[�w���F#�'�%���zit^�D{��߸���</^/:�ϤR\y�������c*��svp��H�Q�J�=��������R��r�&7o;�����S����dO%���8�\����/~64��i�*J���d�?�$�*'�l�~!_{`&;��R� H=2� ��*"���մ�ql��1���ޖ�M�X<�ˮ�'��U�R�4�?��������Aɵ:]�����W� �D�˼7dS+�b�L ��a�?�����߲�I�1�Xy��D�nf;�0�S�����,Q�Γ5�od-,��]��5[����w�7O��ԏ~*6�U����:X�8��S�м,g�pƅ{i!� �0Ku�J�FE���{��g׼8S�Y��(<ΓӾO���.�*� �2C��U���R�gUs�M��'��c�bb�a4ުPl]M���������6,g��i��S���T�~�v��z��wa�<M�m���C��t��r�����3̭�)�N 7�C-�}޸��Y^��c��[[5�כѳ���^*�K����3$+��
��HXVLpF�p%��'-�n�}���B!�e�@L�Q=J:qb��Ҥ���W{^sg	%�?��NΜX��pZ��ۛ��Y:�U�O6����e���*3_���.��hlnG���F��y�4����$I"I�:��|Q��oh^K����_�X�+0���2@s��-���ѐ�6�*�x�Y�h�&�۳I7L�a�W{Dt�o�����FQZy�m������s��v�F�T��DG�c�#���rrؙ0Z�^E7k
��K��H�Y�|�h/�n|~�D@�-R���l��Lu$��<tjt�r��)�d�E���*���:���,U@�  �8J)A�������w`��`D1{��@�٠�I�EV&]7�����k����R��[6L;(<�^�: Pk=w̬�g@�6�°h��*��ʃ��F "�1d��t���1�w�mV�:	A��)�4�.=+M�>lc"ɿ�����<̵Af$�h�R��َ�i��h��,��Vs'��7P����������G���B��'Di��"̒�&�E����\�4�n�vO\�xȖx;W���[B�f��a����	~N������؊�\���Z~qOr��w�v�4���E��}���&*h�Z�jo[ND���=��B�F5�ނW������o�o3�q>h4�|	m���gVR����2v�4NE(2���JJH��8�ua[B��T$&h�Zt@�:B�B��ƪQ��&~��(鮲���Bx�G��DG�Cn�T?�Ӭ΃�.^�Ta޾}���
�"L��d�YW�lP3�'U�3%�@=wM��6�u��Q/Ki�<�x|ڔ��չ���.P���%���Sh�%�W,}݄���rZQ9��QU��E�%�p����< )�/V6;�Z�����������aA��P%��h#f'��(�ڡ�z=������Ã�\�UOލ��1 -p���<��m���o���h�uㅅ#2	?y���*ȋ��ʾ}�d�O�(�I��40>n�q �Isא����������4�;:��a��Ϡ<��ǔ񣨒��F��Z�cm0��"��n
 �'Ț3��� #�f��U"�i�|� �l~�x�n����K<>`��(_v�M)�f���?������v���k��l�t�j�'�g�X���16[����� t�x�̥z�-���ɏ6��O�V��9���KkN#����N|_�ħ����'f堙%������Ds�7BuY�Z�����t����k�*��cxVv^PʚgRΟ���=�����.����r3g��M���W�>&��d*C	�l>M�eq�#����@��O_2%��t��qg��C��2�snP@��(��*�k�:��y��͈��h����Ib`�0%ӚR�/ɡ���<�#H�D�����I�?�e!V��#W�L1�
���LK��?�DiA��j+l�(2�� ��V�_��2QѢy`��ާi}vH�d8�}�X2
�9n?�lu\��ܖ�!b{=�
a��kg�ĕ����$T�%����-BJ� ,b��P��%׾���n)��>8���h�N��ycZ.�����Yț�\����D����0`��0o�mx�֎�D�}�� ��ːsfq��-hᰍ�H��d�e�%��qW��N�&>}����[A�K��<������S���������7h|�#Tz�Gb� ���̦�N�<�D���D�7Gc�҇��-Q=v�K�Zd��|��f����ăl��v3޴ ��s.^��ᜟ7��7�+v����ޥ���XT��YR\�j��ά��!���/{ ������I�A`ڮb��YR�����u��>�/��S�ǘ�x1��5g�6�Τt5Y�̈�N\�B�͊n��7,��*�%'B>F����w�jRS����X`c��8tVZ:���C�͉���v���Zɮ�/p�ي�/"�?I�8��L�O����&���Y�N�udI��~�����\���OIy+���z\ӭ8���єi���69�a,�dp���͡���HtdH���)��`�Y$y�|B|��K�?1��
M6<Z��ˆ�;���[Qb4�(&'D�d�R�ܡ�g�5-����1~	9�g0H�`"�2�^0>6 ��w���B��ΐ�յ��&T��M����	�~;%x��ۂֲ�0�!|��y�©��?*���!����´W�u4Wn�`0 ��!�f��6���Tnkf��P�0p���!w,���[F��d��ތ�;���f碹���Z׋Պ�#��a�V���������M?\��E�����v�����v���C35ܟ��Yn��~��\��I���'m��.���*�d�.bc�ztD��~��\_��n���8Ř\��p��r� j%R%���Z��Q�N�;��Tt��p'Fw(+F��,�`dI�J�^�83��Ro���P<JP:+I�R7ȟ��z�5�6c�	�6,p�8H�rJ�K�lJ��)���#)}&2���ye�MH���Z,O�ڮq7o\.�ߴ�P6/i���!�c��~�*�SldD_�;��Z���H�<� �5�"$��Տc-q��Ѐ\������mX�@���h�' ����Q�4;)�/���FcA$+�]ɲ��Y��Wի�D/ҹ7� �d�b,�U R>��:b�SU孺eI-C�X�����jn��0��Q���W��"L�n���9�d���t�S5�� �	²k�گ;se]T����N:����S��ҋ׽���M!�2�0�ʮE��F�]�c��{�r��7닦�Z���eC<ix�J1��c�����M�՚�R���C���=��Z��"ۈBH���;�|���˴*](WV�P_7R	��D��4��$q S���ϖn~�y&��V�����ȿf���5t�d�r��,�}����*�鐡�>����
���Ӏ)T���o5k05��`����^%%��u#���=+�X�o�OV't,���D�nڷ���˽ a:L��kJ��fbp���6�
��L3sb��w���	��X�;Zc���詔����ʽ6�� �l�U�����<T_��.��l��|�{6TF��Ty^�J�$d>"��:ks|���o'�K�*���X��p0���2�^��?��BC��Y��%뤦k�|h�������7���u]DD��Y�<����Q��-m|���І>���n��T�G��#½"r�~_0�`�3
�)�c�1Y�S]h���� ~rp�@|*������'|[��Tt�$�m
2)aHE��K�E��ҙ���x�,PB�=����_OJ�h �$��,��$�ƽ+1���@C�ҾD��V���fKW���>Ŷ��J��^/L֒U�Y��{͉����§�K�v�8��eY��A��"C���@���D��\m1#�	|�`�D[���M.��8�W}�c=1��|Ԏ�I��e�$�}��M�c��Ѵ�A2F�G��ї����X�3�ϖ�ƫ�1��	l��☳��a�j��E�ld�I$��L��n�+���r�QXK;rk�����fp�ԤZ����w~It�`�͓�K\԰�Z�v/rɯX��T���ǃᐽ�صT��uh�Sj�-2�������MF0-���,РStO�o� k>C?�|D���x��VM����:��q4iȆ2)��J��S�7�M��[=_Ϊ�Oh>��@�r�Brts��������vi�%�<�x]i���G��z�TziO�i�v.Y��af_�}Oo�b
aN�"'tqdŤWYF#3�4�����@��2������,��i�وx����6�C�FPoϗ�@�fv�6� ��,����b�	m��9���U�U�J�v�a�<[܍/�p��Zu�=������~���Z�A���P��:�c\f�B=(�>_���eN���#E�Ls\cFވ�y���-+�P�W{O���Ҥ(��3��T?2d���EvȦOy�9�}Z ��.�(qR�/�>�i �N�s�,��]�s�����K�84lm���Ɠ�*���m�+��88/��P�b��c�^���-
[���UN�rѢ�tyU�}��| *�~���e�ԗ�KW���])�v�]մ��
}���ح���qX�&�]lɼ�j��B��L᣷�������Y�I�/�x���z���-�?��W���YmV�B��n�$��=#���e��N܌����2䕭�f7������D��mB���Z������=��k���`��x�AP厶RI[	��WR��[�.�}W�͏��@5-�8�Wuм&��;de�B����>Hy'q7��B5X[�CX]J2 b�t�MVg��C���o%4P�~B(
��*	e��_y�8����נ�4'�`��4ӵ�/�l���i<ӑ��%���>I�G�e�i��/����
kr�L�k�?7�_<�Sj���(�; 7��%
���#Q'�`]�ޢ�Mv�VE8��i�:�y�����Ip�l�����c!��=~�L����?e���f$T�������B�� ���k8�ڠ񓍣.�)2&�8>�-��HvN�y%*���C��-��7�?����DI���+���y}(�#�񛂢��_�Xג�)ng�P<*ˋ�h�#k��HY�����x`�evxo`�U'��y&����w<[\�W��I�b�^�L$��Ş����b>���-�|��zGٚ��[0������:�?����]j���?��@s�X
U=Q^�ٕK.���f�U��e$�ٴ*3�XV�<�^���)��Ҿ{v�Dm�A��œv?T�QR�7jf�(��ĳ��k{��%�1ˈ��`:T�b@�4xQ�ӡw��P>�2�֮��C&���'g|6���tpl��#T�NW�w�(=�U@�,�S�*oy�B� ��˻w3P
S�yK�p��`� 8��q:0o�^��E����޾��E��p�(��JH�?�t�1L�ݤ|_�&��MY]�u#%Տ�6
�Q�\�/oO�2*+��gz�C8@O.�2(Z����ag�jp����c��+H/T����Nf"�]1T$�d|�x�F@�1ReM����ڶ��6�4ψ�'��}_B*R�Wj#��P��'�i��z9���H+3��-D^�#B �@ ��_��kz����t�a��TF8����	��%˓�����f�e���O�n��]Ri�:��*]����O��5��/�cuȫ� D�~�am�6:s��:�kk�V���IӖ�!���,�5��V�������Qc����>���[���y�&�����������&�2<�?7M��逴��dM�v�����̼nCN_�3l~nn�0���0	W��ڱ�"A�Ֆ�d8�b�֕zO���Af����
�k�"vΘ�&p�>rWx%-�M����Ѝ��N���z��f|�#�w�y-Fٶ���=�ܰJ^�L�9�ŭ��y<e�:��?R�v�_�J�c��C��Сpa�eH4�QJw��G��d������&-��vb��]��\O
�LV:\i��9�"6*��iX3������.v��*݁�l<i{_���;��g�[KH�g@ ���"�[��j��q���-1�����E.X��g���;'�����qI4?V��wf��A�g]��V��l�M���vbDj�*7�_�8b�� 
]�U�8���ƭ�~{Iht�X8
���`n�0dᒣ���">�I��v#dc��扫��%�5������-��ڊ8����A��	�[:`��n����_!��H"!��b0�,��@h'F��N��{�a�ײ�P��|M�Æ<}��E�B���p�z��h�[�p`�m̨��<�ʑ�>��
���	Z���ժF]�;��Ҭ�,,��r;�!���	�S�N��JJ�~g���Ԅ��Y�	�#؃���t���r���X]S�#�8��A$�9���3E��J��D�ڂ�ί5F�~�)�J�*��^ ���Б���w�+�u��Q�V���C��]�n���jUV��%L�J���bKR�qGb��>�s]3�ҧJ��M)X�_�Z�
��o�τ��'�6����Ǳe�{���n_�l�.��l���NF�l�y�
����$.9"���:FC8|�W�o�Y�K���yʗXF�0�ǭ26j���}��Q <ͦ��hU����`7B2rP��D�ל��� Q�m7����d1���I�T%}�G�*�#���r(E�0Е{�D
��S�> �Y3K�he�"櫲~�a�@7G��7��:������`t���h�G)o}EqN��`%#�}�Sy{,�Od�I����#J߯}bW��G�����o��:C1�@����?��V�!�!	V�+6��j������|LqG�Tw��j������,���f�i�f!� O#�<R�"�������;`�mJ�m��	���_����*.������cXgM��u�.�+�4$JI�H�D�����b�=�L�{���1�n[��1�#��;��d�!����^��%�E���~i��W~n �jm�X�;�b��Q�wfK�W�Q���*m~D����>�N�
\�?Zt��r��i����jka�����3�*�G2h���je���ѹZ��x��F+c%�8"�
ʿ!o)�P>jQ|Y��MVH�:#ץ���4�k�2��$J���r;d���[8+Ϊ
�xh��@� B���|�̑8?U�/�߼��g�#x��^G	�� T�����.TM�a� $}
<�!��
�5j"K�d W�W�?n3�a-�靾@��6�}�7�i�}x�����O���~P*���[ z�.����,�|Ȅ�th��9P�Ut����:�?��<|�<���/E��7�Z� �u�d�<��7����A��P[>��^�fݺ/(D �����G��Q"96�\�V�ރ�[�;�-��K�ra��c;��D4�=����{C�2��d�>߅�� |ʴ�y}5��.�(�=�*��>$c� fs7s����-O���܆��4�V��K��Ɇ`W�'���£��rV��w���{B���
����\��(�\J�U؞����� �E$~��6sCF؏]�Kri��I�v��Ѵ��Ee�ӓ��,O��)l�$2jm �hHćϷg��{a`ⴙQ��{x�Rz[�-������؅�Vھ&���8���#�9����N����: A�0��fS	�ۼ�k{D���Bk��Zxy��=T1���0k�D���x�O	P �mRĮ�6�����N�.�Z��(���<��S�SW��&��d����Q�>C!�q�R���ǿvНӊ�2�>Mt��ngQ�C�{����9P��(%��*����ly)��������$�`=b��в�/0���9�< S�z{����IQp�e���JY��B.u
FPUL�y?ҥn7�:j��o(��� R�1L൳q�QG�j`�<�ޝ�Zv���8� �U:3(���ﵫ��l�ij��J1!�/=9��'$�ʺT��E'$���[Ó��QB �R �/؆�I�,��~�o)m�]8�a ��H�Nu���J��a�O�z�&���D�m��&�x��h�Ct���:���3�q�dI"��~@ˆG'yأI5�����{�eQ2��i¬����&�]X�2��[w�k��݆="�ć% ����ѽ���D�|��9z���<+�BǄpq�:���U4P��j��(���=,���Ro貵>f���zf�����3��n^pB0�<��mDv��@��0�N.*T� URR�~jAn��(�Y�%0k{�W�ʌ_����M`U�Gb�d���ʘ���>�U�	g����.�|�g�6)6�5t��b̾��NRr����k���,��3*��5B��-�
dw�U�S�2��˒g`ٗ�8��:�-(����T�W��a.�B����Fpp���e�g??~P�NELI�x�;�&�IYr��u�v�����o5�\��Oy3+�̙zf�8��N�c��R��6�a�7ep�4���v��?�
H�cڻ���Pp�8k_$�}�|x���A�l1i�M�Q������1;���4
	}'83�Z�PRaqM%I��k�h�`���}<9�]�H�%�(�"^�(� l���'`��E\�����(�T�t����	h�u%��$�ɣ�ᖦʼ̳���^�5�*�L�V����Ӑª�$u�X�V�� ���\6��3���,k�ߜ�F�/����Rp,R��Q
s�n]��g.̌.7��5��oB�<���� �1�6��>��Mj��_M�_\黁�����v���L��Ї�7Ci����NnI8���軆孲�}s��Q�dS��bY�mz*�]�3%����/��!�}�7���p�"tr�'r%+��)��(�N�� �
Y�!�>*w�dF����6O�Kkp^��������C�F<��	:!��R�y��Qc&�k��c�ƹ���p8WHO�xJ���"Rw���X�Y�T&(m}��ke�Ñ����O�Ye'��\��1���6%Ai�g9�=�]�����*�k_lw��_Lfm;�R�c� Hn�� �Y2"A��Em�q99��eE�{�{���.Xm�y��b�'�����4z�-�e��A�u�]?TT������.��aJD�>75��Ňb�e ����p��I´�p"I��[Xӂ��׈snw�0Xx��dX��%\�$��X�d�v��I	\>5I �6¨R�e����&�[���:i�@�)���9pҁ���!1��0�ݮ;U$FVV��̍{�p�-�������=@�<���@�n�?�[���щ���M�H�=��n�Z�����Г7����}����]�fq��e�m''����=/����S�կ�p~B�X�+s�H2�'g�~!�tC:tغgr���3K;�^]���4y�ꎨ��f��_�R�	85!Bx�d�w���Q^c�+ >�d�{+�ˇe#V��h�!���nЋ������
�L5f Jxؖb&A�����(PEsXx��-����uX�gZYU�l	��
Z2�&�b6��@�"���6�����_^.�Ll��ı�F�G�yE���
V$�k�"x�:!3�|Co9��K�Vi��/yX�(0��}2����T=��ߐ����!�ah����7��+ɆD%��r8W��QkK�m����cL�ob$��T`��GR�#��0r�++0�G���
�ɽ��Ynb�h ��榄Q~(s�@�ĳ!*u�b���3�`t;Q��c$�)ʹ�E,!�{�(ҏ��.k�,�|sy���J:����bG�x�y�|׊1,��@y8_�:��V7��昋Fˊ�4W۶�F+�H�L��Ou�1(�nQì����2��A��4���dO�73"��{ඕv�7����rm�>�	�>��%֖֐$.N���Z�cs�˿��:�[wq�f*$�4��C}�ٟ.���%�}�т�@��\��ܩʪ��(٫�e�����X���GÒ`եEZ�5������nz�Nm�g��w�;�y��ыf&뤌D���/�~?Թ�e��	+�\
�wZ���ry��'Us���׆
Ҏj@�h�h���j�P�Q;������F&��ޓ7����(�o��">��^|���ԮP�VC}��c��c�w4�.\2�kJ�����F��[3�eh�~�@殦Bh7��W-��s�Π�r��s���H4x�7�)��G�ؚ���T��¬�/X.O��a¦}�(v<J 
W=�"�AUd;)wW�Y13��S�D��@n~	ۥs�b��xiYt�xM:�������P�)�vZ5l���b�,.e��d�c��9��U/Q����'��t�<Ѣ�/�w�NZ+�0����>f�ŧ�u�uAG�P���Y."f8S�(�ef��.�[+ơ��t?\����~&ZB�s-�
뼍g1����Z�"o��9(O�vR+2�z���Y����/�"}(W=M3(����%^K>|� !��s(���S����@M���~4�0����8��,�B�'�.m���ll��sߙX���
vw�����&��?wU�C4�:ݳ `�~��/��f�JC�K���S�Gv���;c���Ι��ܥݜ�Xl��Oj��΂�b���mn�/�v2.��٠�w�x��]z�1�-^kk�@��� K�V�Z��$�|�#���[�N�x�u���t�f��6�&�[D�:�B�>�ZSu%�x�M�sC�k�[�~�x��P׌R?f�7��N<���.�WQƃ����d�n�Wk�^&�kdۊ��?]>>�~q�1��zK�ڟN�$2�;�t6^�g�-�C�y�%�Pq�(@�*�u&��>�yd;	����sU��A>`�*���Z/�����<I������I��eR��e$��\_
!N�L���?m��2w=j<f�(cه m_���ⵎQ���`��ޘF�vYsF8B���p�4�l���	���dlF =���Z!sw�=���B���5d&�D-$ʂO���զ�B[�� ]�}ءhږ��Yb)��8t�j��hRN�������u&��X��z\�<�uDe`�!���A����'	���������D1��.ˁ5��-�^ju��]�n�xe,�d֖�]z	��q�&O�J��s$[�����o~�x1��&��Xi�}����O{t|��z=\���=��}���5���*��h,E�#%�N#A=�:�z��M��f����Շ4�O.?3/��2J1^K�?�Pn����v�~���cu�	T	�R�|�jp�c��m{�����ňz_
`p��b6b��I��Fd�>����d	y����!egr 6�v�t��-�Y�&NM�u�ޒ���D,T�*e��B��ɄQh�wi{bS���&��`��*8�g�:&?�ԙ������G��拮�Cp+& ���?��/ɧ	L�LȤ�6&��Y��xu�6���BJ9�\G�O��+�(zm�8�xS"������_a��SpP���{[��TH��)�51
[J��z$*]|�9�<��1��zMg���2ڬ����\4E�v'�� UX3R�k���z���Y��-N93	Ha8Q�#�^ANz '�=����a1$�ff����T|���.�	��%A+,�,���\��ʗҧK���k�0��*���v�����%|u�	7�e z �Wێ6���I�k������ؖ�#�ԍG$,��L�S��.��"+�I�#�M �JId�Xg�\��ar���K��h�t�5M����n���V%v��Y����B�$C���)��n$�%�K�af�؆�o���8��Hdn.Bbԧz���n(�-?4� H���P���p�b�rMkX%��:�d����r*N�v�e�����zYH�w�v�F�R��P����^|���lS��-�<���:�u�RȂ4���>���c��k�G��p�Hj��JmT��������E&#Wp�,���~���5��O�b��\�I�ou�6 �i�ޅ�`�Ј>lN�*�u�l��%_�R�;��V��9H)g ��"�F�� "�qX���-��vӖ�6oX(����'�66�|�4�쭌 ݥ�(�A5K]�Ե�}U�Cʎfl�D�i7�Is���b=�- �i�����Ĩ��K�XI�6iXnu��4�n�(#0�����W���BV�N�d�z��y�d�y5"��Qkp�#��@�1����2����:�B���F �(}C���,�~��!l�0����6b�F���~{��ר�~�� <�x�I<:濾;Y6�������_��#��S6��	Q�diS�z�N�b30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�)ڜ4{^��C���p�?��|Q=F��|#�@��#(U+�R�,
�ޙ�o�ش`�Lv=Qb8��z�W��+l~���9}�H4<:3ߣpF�|�8�h]��qʵ�t)�H�����sJ��=j��P��
����+�߁˾`�����#��z���5OCP
��z��)�ߎ���m.�1�"ap�G��;d:z�H��]ң�{~L�]B��F�ɧԧ���ܦ�ب�~��C&��aVP�� B�Y��F�g%6��6��oڟL�A�t��Si�#��-[oO\=�9��F� ��&?�mh�u�	^��[8i�Fς�~ޢl��t5C �v�eCh4�ۍıE���YW�y�}���y�5F���^k! 2#z����R3½þ'y�����Hs�a�$��=�|넕P>a��Ԡ�Y��/�=�������Xt�؛ōT��v!|���s&.W��J8US����_�A�����)��{�a� ��O��r�ˤ9UxdD�ePو1�.�e�w��y��M�
���I�#U�j�	J'��S&��=/��̰��r�j��G��+�n8q��<a��]k�/�d*4�_o�{�!�Q	�	�Y��H�<{O�回��>8��}J��{�	\kN�3��E��Zgs`�E�,5��Q�{8�⨣x�~aK𒷍��M�^Xh>�<5g����r�m��� ��B�E��?��V�JnA`+�p�xƵ���f�_k�����H�Z��J�����xx\4�M�%jy� �|���)F�_r ���(�N�qrS�2���"j	Iz/6��l� �)�	_L�Oq�Oy�"��C�5����3K���Lc����:����!��/��X
�9�7�zKP`��\�>�R��\�%���fW�X���}�>��6;I]��AT�Z9=%��ꍱ��	@������o�H�j�qH�����iO�c�PXE-4����<6�QR����ُ漚mb::б~�Ϟ�ԑ}*?Bf�J`�D�q��=��Y}�Ժ�*��;�J��	�fY��K�	�xa��CW���e�a�q���8�h�pD��ZH���)Μ�m�O�N�J?"RO0�������
�c��JR��"_^H^���g�u�覍B���CJ�,�^�Z��t�����;�g�*+l|刹e�k���XA�N�s-t�_���y(�X��ΰ54/�H�Al�W���JDm�,����� 
�<�<�����k+M�Mmh(I=L�PC��$����myu�,���@/6��(��BMw����(H�Â8��c+v~���x��e�ǅF:Ƥ���x��Pu���8xg�K�N�$��3�w���J����u���2�%!�r�`s���Y�jR��ܸz��.�n#0M��6N,��n��Q���ݦ{#�H��-ՃSQ���{6��"��oH9�0g�j���1�%�� X�>մ�ה�R>]��ޞ� ��>���"�c����[}�˻��]N�$"��/%�.)�7�hѸ���C$O�	���h��ORTD~´e)oU7o�.<Y� �܇���W��xa�l�D +��+������mk��3�������V����rj8b5���Z��v�SŁ��̲�v��ϲ��G��)�w�u��p6��=`G���0��'�}��]�� �����ք�R�EK3�`��[�s��7�$Y��RX��8 b�XR�]���r{d���#�m�l�f�؝@��L�?��0��Rye�:�:~��qQ���>VQ��P�C��g��\yl�!���TK2Ų��?�SVbT
t�� �jO1$c!7��`�C��S�m�؄}S�{T�dV�)-^�6nr`�)օ�ē�~�Q$����r�,��-����-�������� ����ͺ�Ĭ�=���kS���h5Rp���E���YJS��`2ᲣT��v�?�K�$����9�rS�n��ϮD��Q�&�⫳ae�2��0���#�٨�n*;�S{�E�A�˟���1i®��(�#@C �O��N&�c��ָ�[����툦LZ����2"f��˕ƑvZ�'Ag�A,fVF*o^7I��x"����v+4�v`ӆ&�|�`�.lo�ftl���V7� ���Ip�
\:�|���!���I8�����)��7G"IG���3���ᚊ�#7$ w��=����v��|@��0�sY�6B�#* Ĩqb<u׎4�����(�>۠�0\3TU������!�P��I��k]���#9�¦����5DΚ�@�/�/X�+�њ��R?���;y�\���;?�״�e�R�)
h�D��4�r6%L�C���}v��U�7�>�Qk�O�ݱ\H�������C��8��C ��1>�&#�[\P���o��㘅�39y�����m�)����e��Ħmj�; ٽ�d�*E!�P��x�?�e��*!5�7���6O��?q��{cz�J�W��3�$w�ۓ�L�5�m�C)?�5}D�N�-Jl�Edk;�ڀ�xL�>��ar����S��XF�К��Q��y^(���&�j��e����!����ߋLLӸ9���W� �x��o���|�:xE�EI��4���p�> ��?%�2��H�F;�Z`ʔ;Ns6�.T0�73��>`�s�ݧ"�q(Z��Z�����ڃl�Y��m洪I����ۧwς�o����>8F|��H+�B;񽴼��YV�F}��%��Lqo����d���\�S��π'[��\�>������ �?a)&h�{�	4Q�[��N��%%����l��5پ�v��4hJJ������G*�Y�G�c���2�5�f�e`����yD����D���P�'O�iԏ�hs���:�=`���
U���a�ҋ���{��Ҫe4����~�nW$��%v7u��yu�<P.ݕJ��wc:HH��q'ę
v��
[]�]�d�ݧ[��T�qh25Ï�H�%�P�hԸ{����ė/�yN��Sb�����+*7z~�V��TEb0Q�o���n%Bw��\�f�*_芏GQ�<���ۢ�:�9�a�LF�w���|L���7S���Q�� �[��)�RQ��A�8��ޒF�?�u�Q�і_��#�ء���R+(D�,&��._"��f�!
�"�8ár�7�+�����}{�N<Q���<�F0�8�"]CJp�
�?)ʮ��J�s�6��<�j�����րu���K�`�#x�Z�����
�C��&6�X����b��1�pp�� ��z
���r�b�ӎ�~���]7X�F^��	���WƊ�Q�ۋ��
����י��0�F�Ʈ+. �XO,Fw������A!���bZ������Y�m����_|�(�3�?t�2�";��I�͟��o�0m�;{2	�?R>ei�GH���3����_�_��)��&�W�mT�uu~�G=ĉL騺�n��اN	!�I	��:T:����N��E�ť�^����a!�f�M��*r�R�
���L�Ѯ�6������[��N����*��s����!�M"���?a�N`_�S��-�q����H��S�b��C�#����/ʧ~<Ҧ����)�Y0B �b����бtE�Zj����ݱWʯ�@���Q2EP@ؿΉ�|Joa!�qya�1�N���-��E�~wʐ`�2!�Ά�Z[�[uڭ��c��Ad���� ���(�ܰG�PBp��b�Y�c�s��˵��t�"C=D�}~�:p�2����d�Y�a=m(�$;����=�G�^ V\�~��{Q���3���/�5�
�{�ԕ$��&E^�@�]F�ie{��x����q9��p$x��@�#��e�ұ{~`��R���ǜU6ɒ�K�B*0�˭[��I.�~�nc/�y�w�s���^� �y�+y��"�P�������1��)D�������4��f�j�g��C6�2�$�� ����j�� w�Q�v�Y�<�� ���2��`���mD@V���ӌ�n(�z�>�>�e�/_��Y���u��0�1E�oGQ2��N���FGK�cY�!��{��+K����3'54�6���5�k��d�j4g@��#��A�3H���Q����	�D�h�ANC�}@�(Ze�����Q1�N��;L{�0lڹ�R��T�=�Vk�m��h�B�����IG׬�V�K��e.~XL���b-U9 �x	�V�s���J��E�����H�e���N�D�����BP���˓��s[���q�O�N��3`�`�T�t�ݨ?lI;��
 PE�孬p�uĘĶ5`�L�ͽ)/:Ӈڙ�V��P����u��:�6�G|<�Fk�O�]�۲ o�bgR�����ô�\us�}?�O���Tœ������6�)q<��x'�\�������ڛ�]��R��_�)(�"n0*t����z?>(j,�ԶF_�� ��ȏoa��5��˷�[(�����U��%��U�y����[��5Z��������j��KB�vݤQt�C���r���=� ��8�fjzl��t�|�4Z����ݿ�o�÷��n�?�:	�zZHZ�����R��0��qi�V�Y�5la.��Էב})��2�7c���{��k3��l�-�
U�QS=0��O�1�x>���WWk�m����e�|��AE��U�j�x���f��
�-Mi��hҥrU�B$E�#�
��8��tS�7��Ȉ����7��?�uQ���Tx,�YML'��$��|q�c߰*�A���N�w/,��IѶl|��)Н�;K�y߈�+��B~>��8˨TJ(�^�l���3��=(k񌙘zQ��3U1��!2���~�-��X�e�%�IA�\T�4��)��c�Z���r�"4��J.:����!��/Ͽr(��}�~H����V�5:�V��4L۷�몇��C����h����ܨL���ka	LT"*�5��9�ǫ&����5��4[O�Z�ax(����Z3�Ks�D�R;*|<��	��xn��5 �X��?{H�e�鈂�;�J����+�=rLUW+:hlV_�Hc�fm�9�Y"9�P��#��*��m���$�y���׭���>pu\#�<b������S-���>MU]����R�\A���e���.)��dW��ko��FU��>�m7��V`�շM����&?�w(����/����V��7;�"-h%���8� ����Q�L��cf(�8+�8zX����}�sf��F=�ҍ�+�;Bqv��e�
 B���ލ}z2uB��O��UNa��W�_O�s�C
��o�������ddR~Յ���W��m\9���P��;=1�
��\�Ed	*	��c��Ú�i��.`Vkn13Mgv�PI��9�ͯ�����#o�w�r�Y�"�W����|���2�t�v��]����q��}&8?��Q=�D��[
O	7*�rS�AS��|�G*D�G��������w��F@�-)rCaz״澄��a#�-�p��x��{�ďW��o�P�@=����Z��3̫[�q(.�^�m=D �&O �Ό2�����α�k��9'Ps�4+t�'�&k�
�eV8�F�W�쇀�[!6l�sjS��	��`���D"M�A�Aj��ݥ4��%Ŋq->Y�*W���DM�{	2I1Е :$�'�ѣ��e&��?͏��Я�T~�4!oU*��'�,�,VIyw�2����/��a�d4� �������׫��������mFq���^�R��{��y;n��!as��}�m����5����� �d�`�,-�'���鵯��������,�>�z^A�ٓAFBJ��#u@��2Ƴz��$�wA���D����MB
9�U4TTf��f3��_v���J��~̔��T�z�� =J;i�z*�ڜ*�HA�#U.���,�mלW"@i�o���c;U��b�C�B-D�����E���V��Y�'�e�P<?�./C&�=���앆�MT�a���^k�P�tu���fAjԟ��p���P���VQ����9�k	Ix͓r����Nt��k$�[I�(�u%����2�]I��و���	�W�&XW�m�U� �fD�u��^�f���>��Ebޣ$�p"���>,ά��^�IC��vpx�������Y�TP�Wf�0P�K��~��W)i��zdƽ(�����݉<J!�����X�A�P|���1J� cWY�VGP�_mN���&��+w��$���k}OlQ����_���dIÖ��R5�m�U9g���0�^li<f�&&�7 �ݝ�JƔ��'��9.�;~��d&�K�(���Ƙ娫���إ�B��� �H��Sd�G��[eMN�$`��ퟞi.�ϥ �6�E�g겪~�g(#z�[^[�(2�ھ��;���+{���4H�?�z���ߎF���>-+��J���~��.Y�S}��τ�%E	X.���4�ub�M3�0z�yN�fy�EqM.ия�/��b�Z��s�K��:{!�h|3��.��mE6@C%'_���x
�)l�{
�� ]���X���J�U%�#�����ۆ��Z�@ty�)r�w���VFUH/3Vu�'uF�&���/�?8���H�נ�G�S�Z|� r}<N�]�>E/�4ƕ#��t\�^�`	r�SʕC�<h-��r7I�*L6��u�{� ��		G�N-���2Q�Z�K �����d�O{�{EB��P�4�˯@��,�`���hn�5�U��������Tc��E��C���E�#:xJۤU+'��%����:��L���D;���Y'i�J#4���\���r�	��Ť�֗Vn֜,�����(��q e2�`���I|6L��9:����s_Y��q�Y;�o�C�^B�pKğ[L0���R㵹<��/��RX�����%�K}UK�)b����@\Z�%�ñfg��Xmp}�j���I*�'��e��gx�%s�,������	(�x���EW�]H��v��f��cUD�=��-�����B&�Q�[�y2�<�W��EX't��V��=D}��Af"�Q�Qt�٣u�"����*]���=�z����f��K�<xx��E���z��٠a�rĳ�<~8�5>���J��U�����D�<�
��m`R0O4��	4�c��? �0�3RE�_K�H^	�gS��s�
�P��,�d˧�yt���M��g�{lI��Ҵ���#�Aʻ����t�Gx��y�s�%K�L�/�,�A;D�D��1�	����'b��Ω�;��j�������:(6_a�ݢ��uu���m��s,Wb��`�6���(|cM0º�V����?�c8���]/��x�r�'�1őϥ��PB#���K�X����e�3j�b�맗�I�Ϣ�`��sq!Vf`�9��Ǐ\j���ܥ��d��nP��M�sD6�����ө�Iw���X{�;���.���܄s�{6����H��gqՐ��Y1�V����%���!�!���]P��>$�+#޵��"���ݖ��Ș4���]�^�"j��/
/�.��v7��)��5f�\XO�O\�Vp���O�Dki�e��7��<&r��I����Zj5݋ҹ�Do7鸭�1�����@�d�/���,TB�V��2�_KVb��I*�i�ʞ�TP��IS�#�����M�4����-��[kp-�=��z��AO�u�o��J�C�.���*!�T�R\3�W���݊$&��:���8#	 /�5R,D��&�dL$�?�D�Z�͒X��g��\񬝲0�'|yD�:D#Ȭ��Q}��>�r�Q���;g���y��K�tKT��n�/S�`�T��o����w:-ѯ�7Z~f`�oKȢS�H'�Q����dc`2-�TnSQ�`���)���6�Q��3�_C��9W-�
d�N�����Z��-*���M�|�YC٦̱!HkQ,����5�С�c�<�Y��9��?��_d��>Mb,l׹�N��DK-�?�Lnk��ϻ�2�No�&.� �N��2���,�ռ�Z�n�&tS�V��M�$���
�iO�=�U"@O[tW��[l����k��B����Z/�~����"��6��s�~Z��OgpUf��o����ۨM"s;.���4�u���|��ߝ���o(Mt9I��Öu �C�I�<
���|�J,!V�v�4�8A֖r>7T"I��䎀�y��w�h�#F��$�F֪k4�>��{%�_�B0{�m���5#W7�>Yuo�O4����.o>(\]0IX4Ur����u!�ꡊ�c�kj7j�Л���rh���<�'�Q�\�`X��z�>��P���x_;�f���e'�{��k��E�)w,h��#�JQtr���
?�j}�vQ#UlH>2|B�\_��	��B`B���TC\��˺���>.n�#��bPy�zo	zK�r�9�l���x���U���ٜ���ek ���+�(�Ͻ>��*rcۉ���	�H�*�be�*�*n�i7�ok6�5O?��Hh��y�W�T���(7NLxB�md�[?2DvУ����R���]��wVL��P��Yf�(����We�=s��7����^u8}�|m�j����GB�ɝ��!�2�Y� ��#�~ �\3��T��k�x�=cE�!��,+���f�DM xS!%{D�;5����Z���;[����ܒX�V��\�� �7�O0('��Z%�ӿӴJl�ug��˴�"�p�j�����<���-�8S݁��U2~O݊�,)��s���cЈ[y\'á,��� +>�?�ױh���	��*[���0�M����l$�5�vv�h^���.���[�YAtR§"w���c5��	���=����#�X�b�<�����F'�ԣ�Ys��N�J=�F����:�/a�9�JID�٘���H�,�N�����>B�vK�)לh�Pa�.q�Z��~:������-�}v��Y[����x-��C�͊q���ã�H��d��L���"��X��ЍT�JCb�I��*K1��?�!bbğ�o��8n�h�w�i��\�*ss���>D<�@��6*P�M�+��ݦw�|��h�K�@+��Q��<���/{�)#>��( ��{ަy�?eLQ&����0#�u��l�+<vv,��M�Bf,á���5&�Z�C8��٠��+Օ��}��}��(<�ɮ�,^F�",8-��]�1R��^)^˦�^]Vsf*��������3���k����`)���n���C����MCY�t��=����f2���w1/(2p{�$xcz���솄a�gr�~��]�p�Fr������kc��0��t
�Ȍ�������F��C+��Xc@w4!u��m�A���vX�L��*t���͈mݱx�mJ��<���S&2����^��FM���m���2�G1?+c >���G\b���
a��ڭ_�aZ��T��[u	�GQ>oL}eO��;�;��!���CTNc��*����X�9�஭��F�Z!!G�fH�D󰷛r5����n��/U��&�Rc�� �%�~HZ�~y�9��������hM6RJfm
�b@.����T�-@I⚡���:`�bՍ�Cd�V��V��F(��E��M�U�=|�0�`�b��t�d�tY�F���X�E�|�7C�sw�F��@l��/=�J@"����a@EN�ӫ-�Y��w^��FQH��J[��k�A�]c���d�����R��(�CG9�5p���.իc	�Q�8�����`tNH�=Xx�~B�Dp�_���ma�q��8�*�4v�=�gN�Vj]��/���T6G� xY/Հ��a{`W$�iLE���T�L�x�iy��ޥ���7�]�8$-!��ԣ|��Dוf�5~t%���0��� 6]�1�_�/B�O���mW�݂M~�U)c�hL�����cm
�@.y������PW���Vnܦ�����d�T��
���h.�j�!H��2�2��u���0X�jH��w�J�vFu�PD� C+�2�
B�E�{DTι�Bmi��;m��넰	E�f���Y��d(D
�D@~1٥>[���$G���Q_G��QY�A���+_c]���3;?J4����#kˣ,��x�'���@�0��f��3\�U��Y����Do0��dCN�S�@�E�e%^��-Ia1NC �O��{%���U Ҳp#�h�W��.��2�h����J���w���K�zL�y�����*<��ɹ90/�x��T��CȂb��˴&�M���\;qeS{N���G�=�Vh&2����+k!�$�$����N~i3���`�@�0i�SWeI���-�W �M�Ðɬ�}qu�Xw���j�a��Q��:�1W�4C����E-4uM�:�M�G�%7F���O#R��o�O��yg�E�)�W\�0�}���O��T�Y����E��@r)�x���\��2T��� ���2�f�f �M)<�0n�<D����z�EG~&!SӶZ.i��V�ȣS8炜�S��_�o�R!U�q$P�(ݍv,���5�Wע|���j&J�K��oݸݘ���'S�����4C�8��j�SV�^"|�������A�Q|���1��Xg	��H��&�R'b9�*�i�@�V�w5 B B��h���1i����c��E��{kG|�lbd���0�]Om��xR����Tk ��0T��� �|h�&E�]چ�p.x�(��a!
��iQ�ҹ�*��u�EƧ�
���/�|xp����\�N�	\Q7G:u䉩�,��,��9M�vy��$jgEq
{����=���ɺ�%,S@�JC� @k�~I���A� y��V>9��˼��J��	Ӏ��}`�Q�Hk�.^��%�ǫ���J�"�Aa�X�R%��u��I��H�f�@�D�w�
w�]r���чD:�6�Gkm�CKFr��N�~��O��%{��:����-<L���>���WH��,����,#�p%����k�	aapX"��n�I]t9c�&���m��H�vOI�^a� ^��3�2�؊�;*C<T���/vӕ�4 �$����H�.��;� ,�=x��Q��L�D�NV�nlHw�%mc���,�r9.E�0龃'l�1h]�V��\"����?2p	}��P��h����O�S�B�&�[���%����2�A!�9��N���J��X� ݃�#����D�m˷WVt�$��"��1��nm�e��C�p����V��;�5h9]����s���Q��p���(l�G�L��Q{�}���ᇰ�z�տ4�B�C�D*8
��w�}���Ba�IO�IN�p�Wڵ7��6
<o�&�
! ���df���W��\�/���O���h1B��\�d(r�	8,���tՙȂ����1G5zv0;��Ǧ�a��͡}Q8:�����H<�6o��v*o��*�u�F4��
�]��8*���Xf&��9Ɩ�=��i�o�i	��rg��S8H�[�u�۶���ܶ����@v>�rW���Hl��p#h����������#� �f�P`A���:Z;~�̿�Oq��?^��=���&E�b���}3�b��kG�����s��tw41&:�g��8��W�#;���u!ʗ5s'�j�œ� �r�M������������97�q��~�*q3�h�M���'��F2���'��Tn���
?aY���@���45��U���'�F�,�wMy��¸`��3����4�\yٰR��'����=�����Je�o2F�x�	�WR���/=q�@����s72����пdZ��}��$'�x-7`�9-ߒ��*�J��Ny�����~Gu�/zr���'��B^��#	bO�Fgz �B���`�b��BL���B)��驥Tz!�*����ܠ�:�ď���� �ᎍ; �#i0�[* �ڜ>�XA�o.�(�w�����W�?�i'�E�m�;i6'��׃C	��D�|���G-1��
)��TN_9�+��#�~Ѩ���u�N�4,�5����>��Q0���UڠW�!�Ċk���8?R�[���/�Ώ�A�ħIXB������zΜ4V;._��0k�0.��Iku܇1)߈Gh*y����Sr���r,���&o��66�1�0����_�*�w��Jk��W0��V�A�_���y=�+w�${��E��l9�5�I}�_���d#���w@��I�9�D�
&�l�^R���0.�wjƮ4�'j'9ȋ�~�a~��������p�Ʋ�~�2W�?����� ��Y�A-��Lɘ�;�eg�$���9`�.Zđ ���E����D}LA�Qz�hg[P�\�tz#�&��'������x�|HtK%z1���8�`�+�T)�*�6u��oG̩�-?F�X��ˡ�Yb����Jx[y���f��E���.�3��١}G&�4��s-A��A;{�ɻ|^=.֖�Ο@��__�Έ��{)��{�۬ 7�@�rz�2�!U�i+�����8G�L�m>�ygW��j�ð�U��c0 �'�,;&ڒ/Z�������G1߭���/��6�<h8�]R��/�c4�7�RA��f�	d��oBy<����Tf����āO����*P�	��ON�A�L�?ZN#��T����zc�iL�{�6���0�ǥ"�𙝣����%�@h�T5��|����.��'��)���������	J�i+�.��,��!X�f"��@藫z�-�J=D���(p\{l;�L��' ���a���Ϝ���5;�(Yv�q�g�2ʻ:�)��Ia�k6怣r���ڍ_��Qq8���I~C܎��>K^>zL
g��l�B�
�hr�/Г~X4'�K��z���\sd6%�fA�X�8�}u�"ꀛ=I�f����<B%L��*W�����q��l�Q��|����O.:İFc/�~W--���/���Q١��i�c�������A�e+}�w��}�avf<�ǫf9�=���w��۝�*�-���
{����f���K��xU-֗j���_a�ѳx�48�=�5��;��������9^�V�P�1qfRʽ��zK���q_����cR��_eE2^w��g����M��$�����,V�ˁ�et���[g�Gpl#�q��%k��EAd��Ϥ6tȵ6��ym�����77�/{LA�T�H�Kr������%�-���]�'�#��S|G>�]��S����lة5��q�jC���R�2+��t}v��qjb�wP�0v�ǿ�� �t2��"�D9sD3���c'�y�魍u/\�I���u�;��Y�[�Ō��1X��g�cӽ�fNGކ#Y�ٿ��n�+�n�)#K3���4��C�B.�ˢSI�W�9���@�ku��;+3�/��$�|�/�Dn�r�aN���@y��e���Ҍ�u1�<��n�;{$���:J�q��F��i����n>h������p��RKTJ��J{��uU%�5a�9O��x�Lf�f�!0��j����uU�e��cN:��Fڅ�5�l�=��m"��D ���ޜ���N&[�3�/`�����j��I*�|���8 #�M��ʬ���u�h˶��@������|:Fޙs"��D��u��>:L�G/��F~��O�(IЮ�v��tg�s�z��2\(b}��O��nT��<��N�����)d�����4\b/��xz�,���0/���;X	h)��n��!�L;zRy���`b|�y%4��1�Ȃ���A3���A��U�Έ����UO���l u�!h_~5m�B�o�]��jE��K��ݗ����&��� �홷���8�lj�W(�]�+|sgI�ħ�������Gļ�E	�L�H�?��R�4���Hi�lV��5?\�a
�g��p��օ�c�Y��a�k��lVK=-,�1�0���O,�x�L�Hgk�{�o���3|g�!E��-��0�x��[�y�
	�i���P���ȑE�Z�
Q�μ��*o�*����(z�7F��h�'���,��NM_@1bÄ$��q)H���!����p��,������o�_(3����F��yV�5Q>��k�[�J;�J��jtԼ#
�pzk����m�����������Ӡ'X�x%嶳��g��'����m�������rj��ƀ!:ܿ'F(�"�Vr{�!EO'~[���>��:�%��i�L�Ê��Y��wQ��ӈ�;�Ό�$����I���a��L"kW��9���&!|�����g�]OH�ak�B��d�3�&��W̿;�}�<����u�Ӕt+ �-`Q��H�C(�9;2a��|�k�p��L��-��V��}H�em�ڋ2\9mXX�O�9�&ssO����,wg�/1��g}(pH�@�o�|g2���S�.i��$eh�ހ�%�A@����s	ɹ��c���U��f�RaFm
`�V��j�����*j-ɧ�*g䎿������"�V'��;�(h ���C�7�Q3;�3�(��f�k�PM�}���.N���?�>�'Bu�롃?�
3V[�vy�}m�B j�O��XNt9�W9���F��
;ro�I�2�r�dw ���W>�9\�i��jl�Νo1�}9�qd��	�����w���J�.�2鮔1&Vv��:������,G;�����2i����J�5/�����F��P�I:b]שo)���&g�e�Z=੪��	
֢r���S7�S�:����-�K��(�H�z�7@��1rv
��G�6����#�-�̴Z�0B��g�W�bIP�P_󈙄�}Z��6�^i4q;�^`�=5 &:�܇a"����T�!��k�"��LNIs%>It�_y&���f��8��WP���ƅ!I�Fs�6Q�WdpŲC�q�M��e�i�(���m�G�$�T{q �[�Ib��g�Mx���x��iMt',$�����!P�?`�U��ҋ�P�4ԋhU=c�'B�,)�:y��\�_p��H´�i4f#��/�PƆ�4�žA���O�I�O�quF�Ө�bR)�(ێ�LE�f�s6���`�����m2��������`�d-���)����.j��_��s���}�z�b��f�zB}�#��%i-z��҇*m����9�M�L�o�B=�k���TY˻��
��c�⽹�<�
&��_D���* Р�i��*�_���A���.x$��
���1W�[oiG��քG;F��u�<Chp�DSڄ�ԛK�vs��l'��bP�s��AG�C������ϕ�ՐTRa!ر#^�I�P��uj��zҁA=�1� �F��+C���$��A���`��Nx��&��c-�9Ҽ^��[��Hc�>%����K��I!`P��8���t�yq���hmۖ�@ur0m^�d�ja��Yϣ�y"2�����ɾh^�C'O&pkZ��?|��l*�Y��j����0#_��i���z�}�`�+��B�ݜ�J�C6���t4��d�Ў J��*WɨIVZ��_��]����qwI�$�Lþ�Dlң��{0_mRkd�ͱ�S� |B9Z"h���tl�9�2d�����pX<�ǌ�'��W9!Ns~Ko�I�^6�k(���9��_��G�{ؘ���-C ��~��%fl\V��Fe�K)$��풴�.ӣ� R��E��ڲV�:��z��h[�����N��n	��f��> �Q��Hm(z/���!������+QAԱ�7��)?���O̢�CX�{X�
k�'��b�
����ya{�f�3Eߟ
.�4�K_աֿ��=s�3�����{��|�).�-��H@6�!_d�Ȉ+x�)�*{}�� 0.�͋j�k@#Uta�T���Kέ#��Zy`�%�����>U;G��"'(�@&���/3l^�{O4�
��Gj�����S^�<O�]��/���4�s�����&	eI����~<����Ν����*���U�c�	���N�����ͅZ_��-f7�̈,���{ئ�C�_����2O�s�#��W�h޴�5wA�S,�݁������Ǭ�>�������9JID+��ս6��3V���B�Ww�������FJV,Q�"o\Ծ��m���L	ŷA;���Μ�E��N,(��q�2C¿��IL6� �����f_��Iq������zCu�p�K7�L�����Hp-���/IlKX�����zK���z��� V\��%s��f���X ��}.*��Y�ZI�5#��`���k%f�-���F������E�D��߲�KQ�	9c�����-��}�r�f֧6Q��ѐ����/Vn�yA�����P�}�rjfU���uٖMTu]֫t2h*pU䳰)E����f��uK)E'x�֗����}�a���Q��8� �NX�t6O�H+�<������mR�n�s�%,��܍#:�v]�XMl��Ij������+���9�(x�
����5�V?��?��A&���eG�1No8�;�B����&�y�Bv������x��O�N{��3�$�`J�P���ǫ2I�����,� �J�7�S���IuL4W��F���4�Ex�:[�ߙ(gJwrm�9$u�\�:�K7G��F��8O��-�c�����g��(�l�K�\� �}���OƫT���'�����)��v� L]\7C2&s�A���.R��1n�<)��n�V*�!T;zǬ�kgG]�Π1��^�3��vjC�߆�S.k�o��FɂUs�D�Z��� '�=�5�&c��)�.�j�$�K�r�,%��'ݯ�GH�wǷ�$8�ljb�R�^|~��|�����������$	�mH�3��f�[R �Ğz�iz+2V#�=5��k��\R��ֺcq���s�k���l����o��`0U�EOa�vxƈx�k�Dd�$4��Q|\�E'�L��*�x\ [��h�
��iE%2�-�L����E:'�
�k���l+a*�\�P��}��7;O���\E� �f,lM��w�$^c�q~�x��y�C֒����,v���>3��t���r�P�y?��6��/A>-�_�0rJ��Z��H��q�ӆ��wky_i�u[���?�mG���ӵJBXs��%:����.~��1�4�h���k�Er'���{�7:1�;���0r��(�~��1�kEo+�:i���zLc��24����l� W�P�g�dYV�Q���
Sa���"��䔽)�9s�)&6�'a����O=U�a t��Q�3`�ٲ̙�;���<H�3�hJ�Ӊ��  ���"H��8��X;G"��1�1���0L�a���GV�HH�,�mW'eڠ8�9"!M��kǃ=��W��J�������#�|�wp�4y��K�\!-�8s�S������G�{E�n �ڞ&A������J�N�q�
I��tᢡm��g6�m�ׇV��X���ɥ��bV����Y:)���&��V|�;
U�h�&���_��&Q����Hk(`1����m�EГ}7��	Cl�Z ճ�B��^�8f�
�S�k!�}�iBU�OYt�N���WNw����I
���o��C~|�����d��	��WS�S\��ɩHr��Ï�1|�6���d���	,�I��KՍ ?��X���,1���v$m8܂U�A��ED���CM�� �Ъfx�j�D3�i!���S����],@&d���&�dv:on=��4��I�	�Z0r��S,QU���*���� �g��=ֿ�t@jf�r˪�<a�3�w#
j�̉�&�_	�|�`��rl��PT�y�T�Z/4��31-q���^q=�h�&���V�@y��V�"k��H����s:�Itkx�&��>[�8*�W�A��k�u!�1s��|�b����f�pMr�b���ɀ��(��6:�4Gq���ڞ��\l�Mo��HX�$��+'AI{�H���v�?U:��X�9����4�lXU�^n'�e,ދy�-K�T�&'3����4;	.٤��ƛh��zP�
�"�>�{6�F�f��}l[R��>ۣ
���؎V�s+{�������B"ĉ��P��.�`�i3-S�f����7�"����H��iwz����pB�;a#������z~���f
�V͏b�F��$B����3T�[�3�8�i�.���.A�O_�X �,pi��K*�ќ��4A	
�.�q��w����8W�Si��G�;�N
����C}�D���)*�kIcC��'
\P����nC�}[�y�Õ��TG\�m^�ՕPx|u�����vA�ʪuY��f��n��G����Z�d����xU\y�^��~Լ�*[�R�8��%���������Ivߞ����ёے�,G�9X���W��+u'~r^Qi��_��ps��>~��6"������~�f^m�pC|p �t��AV�Y[{���]N0�v�9x'��S�����E��5B�5�J��m�8������E�eK!JCW��kVφ]_������}�aw>*�$i����y�l��čwi_���d�Á�Yd����9�h1���fl��n"mA��75�%R��h'��9�Y�~����׊�F���e#�� ��<Ho�-v�Nc i@��o��o����2e�wP$�F��'JT.�� '��Eƣ�2���H�z�M[~��br$������Ծ����f>�H"h�z��<��ьN��+�ԆO<�C���ۼ��W�}���X�0���m�b3�sԸ?y֓�f5�E��$.X��@���ki�����s����o>�{�2�|��8.D�͸�@��T_��i� �|)�<!{�Rt ����d��`տU����:�������z*�,�syz]�����ޟGU�g��A'�+A&��/H�B�0��_
�G_����E����]<���]�ݮ/��4N�n�p���	�˭��o<�"���݌β��r=���X�]	�BAN��aۺNfZ|���Bp;�ձ���{���ش��S$���ۑ��^��dh���5\���H����������R�W���s᫺�Jc61+�_`��̗�h����҇�����a���J��,�Ѹ\i���;2���O�,qT����&��#�(�lmq�#�2x���I��6ԃG�ҭ�Q>_��q&�V���CJ�����KLO�L�����Á�=��VJ�/~i�X��L�K�б
v�G��\�D$%��f�<�X�Q~}��@�n�$I��3�6'��jl%�?%�b���O?� ��ZV�� �f@N@�Ğ�c� c�B�-I����x4��QG����{P��6�B
��M��\��e�}�If��R��~��+�g�SZ�I�j*�>��o�^�@fN�KOxCY*�V��f?,a!���f$y8@����ieS��8��q�e��VG�_�*R�>B�(��zU���aF��>R� �_�@�^�/�g�JX���i�����^,D� �/��td�����g��Gl��<�Z���V�AR?�}�[t6����g����ΥU�/Bg�A�ƃ�����Z�A��qEu��1
��n��ࠁ��"��(��
�e�q8�ڠ>�$mn�|,����"�86d�`(�M�~��qvv��-a�c�����к�����Gƹ��-�P�;��-,&���Y,3�$�sU|��`�*�&ԇ��!�Kv`���OC?j'
0�-�\����n�,qML�6Lv�+H��y�^�{����-e������6��1/WcHnc�g�����A1�y�y���3�թ� �J��]��y��`����ֵ(d�"� �eח�P�h�P��]�2�"��
/�-.>kC7?���~n�8�iOYژ��Kz�$�9D�FCe>��7$Ap<��p��>O�h��� �A5AD�T��@D�ֹ�Z�����bj��-�VaF���8�bJ*��љ���0�H�(�_�9���=χHg��&�>���*�p���=UmP�b�����'��#����5��4�]�+ňR�w3Q
rŐ�ފ�������2�B���p �_�R�ͅ�A�7d�/�������K�ԟ�q��D ��4/�09�
y�W>:̧�lrQ��>
$�8AUg�y����0K�q���znS TX^�|�S���YӇ7��`d��Ӟ�SL����V�pX�d�:�-���n���`b :���v�=�Qb�@���&���->���\������"�mO�ՀE��!��;�9]zk��;B�5g�8g#|K��Y�ܘy2����������9E~����@%n���C��ֺ�&�r���&2�z��Ǩ�.�n�8SYP�v�!�����{`i�����o@�d�0���$ɕ���֍7I�a���	Z�cϹ�1"[�=�����)�Zq�Ag��@fk��o�a�c��"�$��b!�4t��[�-|<��#mo��;t�)��K�� *f%I�Q�
1�|k�B!�*�����%!
�l$7�L�I|_/��vSO����#ΐx$u��2m��p��y�$0���K�f#�>r��w�u���4LJ0��>�X0��%U��� � !뎊>uBk�y��X/��{wr�O��ί��䧦Xb��Ƥ/�Tv;Ns��PSPʻ�i�`ܧUj)�0{hJ%W���r�X�䡉���v�xwU�`�>��>����m���|���<�����W�a�+é>��#��P��o������90ӊ�P�e�b*Ȝ$KCe�Ղ�B�嘰�Ͻ��*������J��{Ӳ`�e&��*��75�6d��?&_��Рp�2�WCϮ
�N��s�L �m�l/?��HD�Q�"W9���p1��U�@L*���v��ް6�2�n���]�:��^����K>j�}�P��Q�/ʋ��n��׫F1 bB0���@�1Ӊxs��E>�m�<�H۫E�/  AO%�/�ä��ZUk�;�2�c���/�NRݞ�p��ק�(���Z�lʿ[_l/q��k��J�����,y���Y���_8��ȁ}��B���1�~Yk�TF2$�%�~SA��oEҁF>Ɵd�S�����k[�4�\�(K���K LX�?66*h9#G	I�3[�G���]��Y�l%_5j�v�h����ˆ��g&Y<i�f���K5��:w��Y���!Ր�������'��{��m�s��"�yX=up6���7a����K�������:3����ϣ$�#D����v,cgם%\�qP.����SX,:17-ÓC����v��[�@����,�03Ѐ�jq}f��D��HಔE5��M���C"ޙ�f��1k����b������p*,�e�)�.�wb�hom?n!�w�m���{�*Tj&���<�s4�w�8��'�aIw��|��\�,��,Q�l�����)��M�����އ�?f�QGD��4*�##�c��OL+�s�,eLC�#P�â���V��kN88��!	;+v�ǰ>��}p�<�`�<F�}�8��4]Xa�ʿ��)�!�?�3sn����?�_ה�%֕�Pߋ*A`��n�Omu�Dt�?#PC�_��y����ߘ�.��1VEp|�e�E��z�G6��*��tz~V8�]��FS/E��v����&P>�b{�
���ea�Ku�Fו�+í�X���wu�>�_F�A6od���������
�m��Ϯ��ɠ��.�T)�2Iz��՗.�¸��.�m�e�2�y�?��b>zc4G���Ȉu~���x_��%�,uzT�@�u���G��L>�cO��<!>��Y]vT�m����L����ծ�YbG�!Bh�f��c���r�����'��-'��X8�S�;�!�|߿>��<E��8��(�ǀK	�MY�gP!Ճ�!�PZ��-��ĚB�#���	b��Ce��&���ӧ���88��x0���b����ekbtz�u/���L���4���D�493'�`@m�P3�JD�ϼ��a�SJNI�Z-�/:1�w_�Չgط�[B�[1�����cYdh��9�S��(/�TGz�ip��~�Xc�2�������%tO�P=y!A~��mp�N���!�m"a����{�5p�=���ˣ���0J���,���/@��?j]{���$�gEs�_�d��`�iZ�¨����!ٲ��$�	��U��j��'�
~UV:��}����h6�Nw��H'B?5��b#̞̋~��0c�&D��%������u��yv�˛��P  ~)�ܧ-���敁��k+�����j�٤ɘ޵2��Gv2K�Q��j�_tww�v�-�G 12�}�F�%Du����ی;9*���y��܄qr��+{�VY��iJ���1Z@��q���;��h�G���Y���P��+��+/�3�:�4E���Nˤ�!���?�@]����)�3����u�Dpm���Nmg@;��e�ˉ��f�1,�0݄{&�(\p��:t�ɿ��k�o�"a7hb�+�ȥ��޻@�^K��_���4��i���9��x�b��kz��=��,i���h���Le�SN���H�o�w!�s��/�������S��[)N���3���`���I������I,�֛�]� �t�/�����u�3D�
Өz�`���i:��n��:����Fu<�g:�=WG�F��O����00d_g�:0&U���o\��=}�OA��Tn�M��G����)���M8�\$��:��n��Ͳy��G�K!��)]��n@�g�zTb�{��;bo��T�����Pq|�q��۫�R��U��Q�!ݮ�,m
�*�x5o���e�L�j *K�}v�ٯq����1g�7÷�= 8oUjozF�_%|�����-�iB���L�:�����	�.H�f��Rh��ċ�qi͝VP�5��E#q�i�0���z���c^Q��Q�k�ml�C+�5��R�0�.O�jx��B�k�����f���k�|i��E�l�?��xI���{��
KviծҚ�_�׭[E���
�9���~���W��._��hp7H�u�r��m�|,YP�Ma���;�$+[q�؂���S��H����,c����B辡¶�?��nyx�!��w��>zK4��J=�u�!'�>h�2�k�*B���M��w�ZSC������X@>%�-���C�i����ج���zrTj��H��:�؟HI��d�7r�r-��~]�V�H�
<Fo:ք���|�L7B�����ò����}��1��پ= �la>0�"�j����9 <�&c�.v�)�OJѦa�q��\33M�Y�YT;��<����Ӗ-� ��Ӵ�HruI靀�;t����5�2ݶL�Wo{�V4F!H؃um�[����9�%�q��(��RlڗS7�����1_[�k�p�=S�1n�i�����SV��<�j*������$/A�ـ�����p؊W���a���X򎔓m���VUR=�����R���h��pE�bi���k�[��V�a<;��hZ���%����Q�q�u��(-.#�-O�R4�}�䄾V�)�G ��@��B�t$��(
��xB�}�8B�{1OF'Nv�W{HL�ȴ�
�Ŀo���+���u�d�Zͅ��W���\�G���_���*K1)���1mdd��	�8��5vt�Zy��bq��1hR�vq�7�����)ng4�ɾlk+�6��W~﷜��Y������
���X]��7+��ɗ1&��l'"6=��l	�´rH:#S9���|^��^���*�.���@7K�r8)��I����|�#W�T�v���2�迩�1���^�\Pa���~�Z|�M� �/q=|^G*�=�G�&�`χc�Ù� kޣ{�k{��N��sg*�t8Ԍ&`�Rh{�8�Wһ�X\ !KD4s�D���:��t�քs$M4~��M�v)�I�xڄUq��{��лii�M��"�E��O��'nv������:0?b�/���)\�4��U?W�'C�`,��oylw1�a9�ԋs�6c�4(A��1�e��O�G�w�=�K��X�FF���jAnR+C����
��m��69s8lX��,�\"%�/���w���`X0�-�aS�+n5��Y��]���5ֶ���z_����B?��#
~1�g��za���^��D���5dV�B��ԧ�6`T�:-�kbJ�%�l����Lf:���oO7 ��iQrO*aF���4A���.�� f2��b�cW���iH�!�X�Y;��S�w�CC���D��\��8%�x����'Wp�Pw���C-RC�L��FE%�{�TTx���^@)/Pe�?u21⼚A��F�����܀�|�����`K��V��Y_º�R4,��ٵi��O��M��{-5��9���uFʤ+�ndfR�ƨ���Rz���;�s�3��o[��8?�3{���>���G`��0-�*�W��s���M��9��z�z���l�BC�U#���k�z�~�����g����G?�0B�n�n�DT�ܟ��D�)	�?��Pjv�e<�sd� VǆiU�5*�?����LA��.�N����f~�W(��iL$ ��
�;Όd���kC���DY�����c������y'�)P{ #�ǌ�Cߜ��ʕ8�uT���[K^��Pi�u�Շ���HAC[Ԫ��5�����n�⯜}�Y��kNX�$B8x��H��ϐg����[��)�^%,�9����ʎI�1.�6Cj�BЈ�5��\=��J���ux�`^G��C�!G�_����"��ƫ�_y�ϻ�^ެ�C���p��9�E�߸2;�Yl���C�0)���m	�p����"��k�{�"9{Jڃ����.�j��'Յ��J�!NW���V�__&������A�w���$�����l�杍�c_�^�d"�������j�9����r�l�:�3�$���v�3ƍ(|')�	9g�g~Q�^ݍ���� ^�s&Ƒa ���$��0��!% Zk���3��g���BeF�b$y�.��%�.�=P p�E��c��@�z}�X[6v�oh���n���
��l�Ǘ+YHs��z���ߧ\ƌ�X+W���w���T�`�K�̨	�e�XGݬ�m�b��ԩ�y� f2d�E��.��k��W�ɢ�I�s��C�L.{��|��.���^g�@|y_j}|��P�)�4{��� 6�*�Q�C��6U^IݖҎ������:]��yfҗ�pEh�oPyU�����'�^�&�/yZ>����M~G�d@�T)�Y(�<�Y�]��/�X�4��I��
J�w;	�����B�<�5�q��㸤�é��t���sf	Bh`N��e۫��Z��s���1�H�B{^�����R�$A(�����g��D�h�-5ͦ���T~�S��=
��j}h#��KL���KJ�ޔ+@9�^U��9^j��K|�ݘ{���� �hJ(����c\Ě��i���b�=�(?����s(%[qX�2I\��V
I��M6?�������_r��q�p/���C;(��	4K}��L	x��K�"��VyWj/O+Xp�b�]��K6
C�������\2 �%�,wf� eX�4}�	��f�I���%��'�%�� �3�
�)�����L���:����g��O��c�f$�b�-Z|��X*��mQ���(:�u������J���2���X}�=�f��j>��܂^{;'�:��*�����T��-�f�Z K�x�+L��~G�W�a2*Ƴ��8�7�P���&y��,t�B���p�p��R�d�y�n��0$�i!iR���_�E^�ҟg�Op�L���i�O,�
� ��tU���6�gҊfl"B0�ˬ���JA�cN��t'��v��_ ��&��-�/�,kAR>���e|�?ϒR	-�Y���7΢�a��s��Q���8 (�}��v��is��@�m�x\,3ia�ӵd65�(��M������Y`����JcQ�������x��������^�RPm����D�q�͔
O3Â��dM����[^��؆!O��`�fԩ `7j��+��΁���n	:�M�OW6�i����7C��/�{��Y׃9���Lg�6�Ǎ�#?H��gnڗ�vNi1+z���66�h���h��f�]�hW���L�� �9�o"��'��͝���-��_�]4ӂ"Ö�/��N.O�7p�P�Y5j�W�O�_������D�8eO��7Us<�:��B�����Nn���n�D����Q�?�����W�]sT��;��1~V2�<���b[\n��B+��
����\�B�X����O��[�~p�PT=ƒ���Ů�j���;�Ff�e`��|A0RU�3����A2Q�}�o���0�Csğ�) �QR%���Ҷ�d��|�|���5��+M~��is�������0��yK b:�f��]�"Q:q><�^*ߨ��g�� yR�?��0-K�k���<S<:�T����* ��
��7�S.`U���W�S}ˋ�*�����vd|�-D�=n�o�`S����,�nb�Q��m�XA��RɄ-�jI�o�;��o��Z�&D��@h+�h��Bk��3��5x����%�q�Yy��
>�֢�F�����J���qf���ndo��Ը�J*&��k��/�2$�L���¼!$n���S�7E�'R��}kr�l�i�^��[@���m��t8�I��^?��R���IZ襝�Y7�"�H�3�V��ZZB�g�f|�WoD�#�ʤ"l�i���4����,T�| �4]ko�zt4J���V �H�IV��
��|\��!���/Қ�v�j֏��7m0{I-��ٷ�g�ؚ��i#�V{$Ɠ�֣��!Uu����0�g��\�h#����9uh�84�/���Q�>��.0�-7UC��ʃ!p�r��M�k�`��	�1�LFg�@6���R�Q�X����7^��+�?���;�)�A0a:ךէ���)p˽h���dr�<�O���`v�c:UE��>+!i�u���B�u���v��������|��>'�p#ވP��jobq9���=9A����������g���6�e�3��d����O*+q\��j`��C�CM�e�l?*�d%7$�6uy?W�7�!�9�r1�WԼ"�}@��	�L�_]m��?đtDO'���7��k�f!��&��Loa񇯇���C��w2�6�W�Q�f�^Μ��\�jг��������'�rr��.�|�� S�����
�bƍx��>E���������;� �#%~��8��+CZ��~;t%a�K���
ӟ?����C��ݿ( ��Z�j��R�l�֩T�Z����	���]O���i�&�b8l�0�..B�P�"�Y|��Fc�u%2ܞ��Po��i�����pkS�v���'6[�L�\9G~���B�� � �?{h*ܳ	Z�7[� [�Bt���"�l�Vb5�S�v�(�h����#��-�YS܍�����5�"v��2��S.�I*Z�N��9��'u�=�u��s��I�US=�f�g��L،a*���$�C����N���~x�T�N�P��v����.!Y�"��.�߸�D��:B�o��!8�?�DvQ[�=�J�rh�q�Lq�C��u,$H1��D��ޯ���ѕ�jmX�ߑ���*�b׬�)s*�Ǭ%N�ߓ<b�l�o�-{n2�Vw�.�c�*�;K�m�<{e��H鵄�8I�r�xw�N�|��ɝ���Q��v��Y��N�)�{W���&����?��YQ�w���d#{Ţ���+,�vޔ�|�3��a�lVL8)J��2�^+��g��{]}��<wd���F���8X]i�]���)p�咰ms�rm>s�i�ׅ�֦�R߼�`;F~���r��y�����Ck����_������G�1�NWp��zkz�6��؃u��[~��]�&F���/~f�=�a����S��
+$�����%�FHP�+T��X5��wFb�P��AGXn�H�d^>��|0Ƥm���}|���7�e�$2z&}�&ʗ�35gە8Vmj�H2�lY?}*M>�NhG.FH��hY�+��_���֙���PT��;u�)�G#�2L����ԍ���!����*�gT������7�����K)'��x���9!�'�fZ�!�rǉ����w��c}�kYU�����҆�ߐ5��ߩ�'��Y��� EM�:��_��4�j���`-�4[�s���Lx�b'�aC�	��׿�����8e��)����0�jWb?p��|pt+BF \��=��צ�������s��
@�1��J���Ta�F�NzG]-*|���w��N�^S�,~�["jm�ӂ�c�wd��_�����-(���GKpp����c��D�Jbֵ�ht���=*��~Tkqp�Lʕ�Iݥ[a�5Fʊ�ƆN=��J`
��|%��Ja#~�f�J�R��/�WJ��s[{r�?$��E�w�&��� �i�dg�1������D�e�Ɍ�=�6Y� =F	|��r8�S)K��l'.�r�����ׄ@'*(r(�X�9n��5�#G��fs �"=7��XJ��ȍ�	PQ$��'}Zl{*�`�q-�I^7�G=��&��m�S6�ݙ$ޓ2�kk�|�>�sW�[t(��&P_wX�[8���W�b߀H�!;g�s�����ٯ�d9q�c:M���۫)�f���9����uqr����ѻYt�M�v���}5��?��'^�� w�ӗ�?R�Q���U�Ӌ4�\�U/Jp'3�,�J>y\�͸Q$���V�&�94���!�gƸ�"�7|�g)�;�ӑ�F6)��Zv�R���2ܾT���c1s(7V��B�Li���ĉ�9d�	�`Ho�-�~a�)��r��M*�%�i欟zp[��D?B/�#�(ǵW��zQȇ�������Tu$B�ާ�ѩT�3��[yf�������<Wj�ћ��_<' �iA[�*Q ��1A�0^.�g�V1��R�)W�)bi8�ҮH�%;����gR�C���D��*����h���'GW�Pgf�3��C���6$��k��TD�
b�^0 kPU}�u���KUA��t��q݋
	�u�@�-M�����שM��x��z���Op��p@[W�_%%������8�w\NI���� X�.[2���wRu�Z����u��^�� �\>��,�ţ��."$B���^�;�<^���Cۑp�d����u��Y�	�����0��;���t��؄���Ƃ�����&ݎ��J�(���=����}��_JV�OW{+VLo(_�@��v�gw;	`$W'�0�l��_��%__�[od�,S���~��O�9�t���bl�8@��?���������y<'�(�9S�\~�Y�ɷ�P�)�U0"fC�}�۫9.H����i F����F����cl�e2�$�پ��<p.E2� �E���O���eKziA�[{�^���c� OҿrU�0آǃ�H��\z�&����-+�8T�cw�������O,���
UJX��
�YG:bp��ԕ�(yS�?f�EQ�.���=�f��p��zsx؞���{�_�|x�q.���ʬG@hl_���ݮ�)q�t{�L= �?��=Z��]v�UJhS�w�Ȉ����Ig�y�$�\�,����Um ;��'�O&���/e;n��>�*G\�e�@���|�<�;�]�/�eN4{��I��0�	�s��ZC<�%��w<C���p�/ �`,{�U�	.77N�yۗޫZ����_k$�>4��43,{����u��ǐ�D���e�t�0o1hP�W5�"�EN�?=��B~�r�q�穂���h��J��+��1�J����"��	*�Iᗶ��l�J���ڰ\C��7xP�r�5ũ���<t�q9�� �A(�"�qD��2�_�tlnIX46��~R��{��_�4mq�G?�4� C'j��u��KiDLu���7H��:�L�Y�/�l)X\*-   ^   Ĵ���	��Z �vi��:'��(3��H��R�
O�ظ2a$?�K&����4`��̏;Y�����,�P���#j��6��¦�޴J�������'��Ɲ����dL�KOZ��P*~�n��ѥ[�$K8O����7;�b�O�I� [�8IH����5�D5��I�=^�;�M�LyR��	�Ay���0��	D�+�t�т�/���`옅a��W�o*X��p$�j���Ċ�<j���^}b��"e��2d+!�ĕ(ǂ�1mȮ&�"��xrd0hK�yZD��tf@8=���2�'�9c��9E�8tp��с\
��O��"�(O���N>��&�8� t�d]��P�D��<��=��"<1�AD-0l��u�$FgN�i���j]�`���4L��I�V� ��P�W�\%��Ɓ"hi��'QjEEx�/�R��� ������=&�ć��1m�%��(�t��3%h�A���4��b��Ƞ@O�U��%5�	�bj������D��R$kx���ʲN��a�j�<i��5C-�㟰l�]���#�>�F�8wA�p>�t���	�n��,�|T�$XG��/$�4���'���DxrKc�I4/�t²*I?��\Q��*2r�ɩU���9E�Ʉ ��Y��"P��˦&B)nN2�Ę%n.���NS��3�a(�]�Jis0�.а���	n���E�L!^�l�+#Q���&o�0�H�Od�����?��'��D���L�(=f����t�8�g0��,zJ>yw�\���T�<��퇱 B��D� &@ܼ��%K�7�P��'�ղ@ ��G�!�$k� �  �                                                                                                                                                                                                                                                                                                                                                                                                                                      �    R  �  �  &&  x'   Ĵ���	����Z�/C�'ll\�0�|r�'a�	�Dط8��0b�
�<�}#�'�t4��B�h�dt,�:?������i"x�	�-��K����1Bʚ�HH�� Ҕz�J�[�.�0�|)`��u䨉:�Œ�_2Ii�$]�-��s�	��	-�i�V���LX��92��6�x)����sA�)(E&X�9צ��
����q�`˯do���ЂL99}�4y2�E�C����>��(J�"���U�i�����m�<�e���Vk�$�r���3�,���E^�<�Ѝ3?�0���x"���,�]�<�BcQ�P�nЈ�"R�	cT����M�<YDc�r��1��Y�����F�<Q�ձP�҅����*
8�P{6�B�<鲆
(z8���J�%~A�C�N_�<1�!+��|�p!O!gƖkB�F�<��o	�;��B��[;Q�xYq��~�<�և�+}xe薋���b��d�Qf�<�!��.0� �a�=5l���
d�<��"Ι%yMX$(��^W$���|�<I$l[?E~*�l�!Ha�T�C�y4xF~8i�bL�qȂp���y�)�	{O�|���
�txf���J�ym �}Y�*#*��7\�@V$C7�y�M+,:Ѐ�JB�9�0C�gN�y(�q�:�$�M⧄VG!�T'!w���3�X,B���]!�LJ�.h�wD	�6�a�P��(v(!�D4 ���H�o"ʁY��ѻt�!�$!W[V��1΀! 1��F_Z�!��T�Ms�@�/��j���wFòk�!��D��(��&o��B�/E�!��q�%��O�2�&yz�΅�k�!�D��6��<	o�R�(�`�M�<!�ĜRq���Wc&V��K�-<!��yy�����b$�Њ�t/!��H�fؠ���0�����V9!�C�p}܈r�j��Se<���Α�B䉭W����KD��	 �3|pC�"Oh�q[�	 �j�h]j5�փO-�C�I�"�� �S������0��C䉴([4��BH
C��]�2���1˨C�I�3��c0�N�j��q��&����C�ɸ���[2��1-�Q&�̧:�bB�I.t*�]�7+W(8C�[�/Р"�2B�I�r�@�D ���H2���
B�UCL�⋀2:*�b�;|�C�IRU@��m�	8���k��M�BB�	/���ck�u���"D��!:�C�	8W%����o c~�E�D�î�C��
=�x�0�E��-"0�ˆ��7D�fB�	�+���ħ�bm�V�D�y�hB�I;=���+� >�@�1/�4+%XB�	�~0��ԧ�3[i.i�0(��sxB�I,\ ���d�ѵ3!b���S�BB��9�0H��� C'��Bh��)�C�I\���ao� �Ď���C�	;A�d5`���/}����C�(%�C�ɯmh|dZpe��o��0��-�eA�C�	��f����N�h�\�'F�B��C�ɣ;���{LG�s�r�
fσ�l(hB�I�v!��đ$8)F��� �Ju8B�ɣ�dX�g$�6%"��P�S�&Z�C�	��PE�e3}�]�g"ݯ~��C�I>�a��"�1zr6���"X3ZB�I!^0���"#�-<����DX�L�B䉛jwL��JݳM]�X%��`8nC�)� RL�6g\�F�
��f�%Z�"OmQ�2����w	I.80��"O����,���"��c�N�3"O�U��M�B��L�sȞ�M_r���"O��V�>n�A�l&X]+q"Ox In�>�j���	��v�lA@"O��Ct��C�����4E�f�+E"O��1�ED/Cb4�����`)1�"O(� ��bR�@��0���1"O��1BոL�|<"<H�Hq� "O�k��&S<EQ��-���%"O� AqВZ�RP�%����S�"O���cLa6���\Ȉc"OJ0� &Q�z��@I��[�_|��"O��V���:C�t��GB�U�p�i�"Oͨ�k�7���s'��1�U[a"Ov�+v-N3�j@��e�[ߚl� "OZ�b/2�tC1�M�dȞE�r"O8��O�#3�)YE�R5`|�e"Op�ʖA���8�f	�}���"OB�xT�L�P�a��7�%!�"O�8ش��)��t��닦,c�}�3"O�)��M͜�� ��JկZ]�3"O(���	�*�\XtI�xJx��s"O�Y[&�K�AT%���E����"O�-��-Q0 ���K@Kۨ\{XS�"ON9�F�'Tࢯʿ;Q$��"O|Uc؋e$�r� � V��}��"OHp�)��.�a�
�%O�� "OH���DG
�B4�q�L?D�<�*�"OJ���
.q�u
�9�>�s"O�K�%\,NHw	ή8����"O6�˗�SfT����/
��h��"OR5�A,!L2��OS1s��3D"O>q�&I�D2��bNح)���%"O��F��1&ʄ�#��t�#q"OX�����IZP�����3�X��"O^�U��ZrΔ��D���"OL�auGH�|�P+�Ů���"O
���Z3R����鑘b%Ъ�"O���*��? �	�hcܬ��"O�{U�;ø$�ceH�e.���"O�)��ٵj�����Q3'V�@�6"O��Ң$B�O��X�j�ܑ�S"O�Ds���4��R�hN�C��D�G"O��U�O
.1���SD�2��"O�$�R�?OH$q6/ҹ~0H0��"O"�SGF\=RY�#�A&�;�"O,hRe��9Lv�]�%�������"O\�s�M�W��	1��)�BP:'"O
y��D��-$�S�0e��Xxc"O��"�'I�pZ~=2�N�:�6(�e"O�1�7Y�i�PO��85����"O�)��͂&�ikw͕9#�2	�r"O���@�R�������'�,�i�"O8ɱa�٣g��U(sA@�t��e��"O2��SƐ(/9�]ЕG��I� 4�"O ��5������&K�h��\�v"OdiD��"y:�3�>*�"O\�K1�H�]
���
:<�P �"O��X��3�f!CvkFq�d[�"OD������RA^��ֈ$�"O������B���sf�G䨚�"O���Q�Y�8�
�{`�϶X1��ڀ"O� <�G�S/N��0��3M�,�R"O�T%*��x�V!z���|��"O�$r�)��=�l�j���
0�2L�A"O8���I�hV��  ���0�.�c"OT9rn��.�{h��e����"Oe�&o�$t*8Y1�9b��"�"Ot���6���b���bVb�XG*Of���̌����h�H��m����'9:ٚ���-�T� ���P���'�hiC�����K�^0�	 �'�>�bH��^�։8`���R�v=��'��5C���t� �:�ڶi�'��@feC,Sf�P���6F� ԋ�'�t�jb凌0��=Yu��Ky��
�'�pB����<4�$	�,O�Y �'P��c�a�7u�,��ۋ
!F��'Z.@3拌5gf%xg/ܟ h1��'�}y�)Z�=$!r�E�A�4�p�'��xx��o�& ���(w���0	�'ђ]yA`�)"N��"���Z�Ν
�'Q�������!��O�_�* ��'����a&N�{���ѷBR�<�'�@�0�c��,#PQ�4,̋L�x=�'�(J ̊�.�@[�`��~X�`	�'�d=`2��R	�mkƃ��w�+�'��� 針ϊ��1�OOTC�'�6�pED[�.�bp�ƌ�X2]�
�'� Yi�%;
*��E�/_k���'�hu�Ǭ	!f��,��a�G��\�
�'Z�T��x���U��͉�'H��#����xИ$�U_	L� �'�z J�*�&j7�ˤ@�6W��;	�' 
u�E��& ����"Ҍ]	z-��'TDQ{�!��_ H��9b�8�'�Xbc	4qw����!�Ϩ��'� �CmK�o�`��g����A��'��)(Eg?z��-�!˻5��mQ�'�<��Gˋ�[�H`��З7'�t�	�'��Hr��33Z�J�a�>#���P
�'@|	H�i2yN�@b@��1�	
�'�B��e�{�vlx������'�a�v!�+�Is�̝�Y
�'��djG� }��Y��K��3�'�v)�!i� 0��́r��$t��	�'L2���B��(�`'� � �"�'ir@�*M<nh��+Q��F` �'�nL�A')���ĉH?����'�d�`�"˘?+�� �h��<���
�'��q0��Ǣ\f���7���3Ϭ`�
�'�f�[���(U��`����#�$[
�'(̪�E�.\ԡ�1
L���j�'~E�s(*�ԋ���O�f���'��yp N�%f�ơ8$�ͧo�`"�'�49�i_���E䋘�8)����']�u{�l� �*�ɠ�3>1��'c4 v��@�T�JC�:�X�B�'� ��K�/��)�s�*9�\�	�'�$�
E`��1�tAYC��(t�	�'�0�j�D#H�<�ӌ/)��tY	�'4�C,O�=�<�g+׊5/���'4)ˁ��,։H��5�`���'X�4���X
G���iB*�o����'>��r�֊.���u����5!�'�A�(ON����NJˤ�+��� ��H��"4	�	۸rb��t"O9iE^�U<Mp֯ϲ=��� `"O�\�v ��0��E�3��\�"80�"OVI�
[�8p6MYG*�<X���"O�a#�+�o�H���F��Q"O+M��l4́1fO��{��W��!���:B���H�"A�ls��ޮ�!��T��*1�	D(y�(e�!���7 ������ß"c(���ʝ�;�L|�Z�����	�U���A0f��M���z�AS5}߈C�ɨ_��y��$��諤�;GO�B�I`�l�s@�"i��C��B�Ɉc]NL	�Y<,p>��B͍!_ B�I�"(����;�J�*ׯʈt��C�I�'q0҇KL�k�Dl�%���7%�C�ɘa6x(f-T��!I�R�JTB�	�no����N<J_ar�D��$)�C�I�~��D��A�$9X�H�3:�(C䉛62l�����:Qs���2A]t8C��
�QČ�uH�m�����4C�ɰ4,�9��/�}�DS��8HC�I:s*�$sB��}��M��	۬<XB��	) l�
�ϗ <TԽʁ�ܝ�\C�ɰw�,02��"M�dq-�#qC�I%A�4��2��=���a��U�[l2C�	kS�"ң?D�9�%�&V�C��#W�
e�aS=)R`�	`�`,(C��
����c�@9H7�1��+�L��B�	�7�V4��KD%���₢͇*��B��pT\���7bJIR5Ν,U��B�ɃG��8�3�WvP�ȳǫ�u�ZC��C�va�pIW6IfX�Y��G���B�ɯ�
���N�:J2&Ѐo�r\�B�I�Y�d����<#d��$�8D�\C䉾7ܴLRG�§:MrӧN�q)^C�I�>e �b,ؘld���a9U�B�I1>�,��<��T�eFL��~B�	��ؘd��l����i˅�xB�ɯwc``BƊ�9j�p�� ��>��C�2do�X�B���d4�u�˙nK*B��#Q��E�E�V�A)<*��\�g�(B䉁R��� iؿ6�+fě4B�B�$\�� ���҃B����M3�C�	L�f�2v!˙{+*����6{&�C��'^������U>Č:a�ȵ{
�C�ɹy`Jpɒ��	d׆��0��2x�C�2w@v�CƬ�-�\�+�f��D��C�0b��a��ϑ4���`�	y/�C��h��b�A9`���;ׂ_&"�LB�ɖ`���p��^33<xu㥍><�&B�	��Eb�J.z�H��h	�y��C�)2�H��L�Go�Q��JC
M�C��<C����E��N ���l��C�	�\<N��#�G�9�n�!���[��C��2w@L\9p'�!&n:�t@�t�C�ɸ�0���H� �5�h ��"O�1i��$a1�%��N#���w"O��။�=�;�N�dnI��"O4��1cM�{jY;��@�~4�[�"O����+U2�>Ds�,1�(�D"O�,��d,
� �LU�e�h��"Or�X7��'�Th�����Ф�e"O��
��ݫ*|�!�*_�{p��"OV���mځ-(Ah���fĭ9�"O� ��Au��!pe�r�#VmC�m�"O��B&D��qQd#)�졐P"O>�&���T�
	�b^t��E	�"O�������l��YG�&���"Ovѓ1IZ�~�B���<���"Or\�Ԉ��Q8��Ǌ!;�"�Ѓ"OL��"A��^�|���}�̴��"O�(��*ٵ5Ȳ]���="1�5"O���#Ip�Q2��E�1�"O�Yk�d��CtCƣ�tzd"O�B���:�d��vǏ��~�"O^�h��!�0�r�EQA�|ZT"O�e�b�Z�E�X�7ś�0�v�;�"O���קÇ ���c4��3	nd�H2"OA���D:]�:�+�dC�WevВ�"O��鐀љS�&�1vAD�j>pd�w"O�Ѱ7O����V�X#���%"O�|�$j�{[`��$��K�80�'"O��c4&ǆuw��'B� j����"ON=�/B�H�ോb� M�1[g"Or�
e���ޕzf���5�
ŨT"O���g ���}�a��6���[�"OB�Z>]����ɋo&lA5"O��2�.ɥ"��E�'��8&�H"O
�O�!|1�$���5W�8S�"O���皅t��p!	K�����"O�(���L}����+D��}h�"Oj`"��
�4YR�VO�"J��"OF]�f'J�~{���Q��-j��"O �#$jJ�& �1t,D�o_��(�"O�$��Z� �:�+��$<:�S"O��Z��7"M �2�X����"O�0rfhR;j��T FfE,�� pt"O<Ձq�٣<a��Җe��|��)8�"O�Q`i��~�˳N�M��E��"O�X��]!j�z�ʲg�$���"O�RQ���:x@�&旯Mΐ�%"Oh83���u���@��1r�b�+�"OBU�&e	�Wr�c5��rߊ%�d"O�[V%�	�00���NΞQ�"O�Ѳ3o[a�D��?mZ�*f"O$�V��/?j�A5BO�gNr�a�"O�Uk�e�xz��O�6C�I#�"O�����״��狊�ba)�q"O�����r8�r��5X����"O����Ώ�*dX�RIƀ@T��`1"O@R�+cq~Sw�֨_>�i�"O�ɘ D	T@��� ̯Tŀ�		�'�J8�Fo_;iQ��HS
�b9�'A*���+�
Z*�S� ��>�+�'�:�u�
~j���rg��	ޤ�'�"�b��$KU,t@��M3���'��8�H��dK��Q1�^~
@��'�hh��Ȃ���yc�ȶ�nL��'�(���8�ԅkU��x���K�'�P8��
LAk���.��h��`!�'��j��^+q����dgN^�4�8�'`�A���{��e񠝉P��h�'=b����b��%
Q�]�LRFD��'���Z&�@G(TK���G� �
�'�|�����<�8� #�P�r���'���5� [�p�oQ
	?Ҩ��'��iD�������E��t��'���hAe�0{A�]�@!��s�"O� ��it�̮w�X#��U�i���p'"O<���F]�h�H����E�)�
#�"O�H2�� &�~ŃW%I�i��8��"Oּ�Q~AZ��A]��M{�"O2`����;�e���<?v&��"Oq@
,0�H���9���r#"Op���h�R��%͜A�X�4"O�bdm��.�n :��¥w|N	sa"Oȅ����~8ȡA1��q�A��"O��S�R�@Ъ�����! X��I�"O�u� �0f�Z=�ꗆe�
pb"O���G&ɶc;���J��t��<��"O�Q�ggd\��(ң=�zm�"OL1���>V���Є�D�bΦpa"O�lS�m��?����W�`�
��"OPy��7	r,P���"�xʆ"O`�������X�=��Y��"OT�ڥ"�*\xi�� g{�,+c"OP�Pq�C�F.6�Z'��^���i'"O�����<O��Ex&�Z�Cy(U˅"O������z��鳒�!<O`�Q"ON���O'Fp����Ȥ[6�-XP"OJ0ˁb�>(��ظE)��T��U��"O�Ȁ�+��*�*%ZI��w���R"O�	
���R��D������c�"O���!ڸ��q*�ǋ�`����"O�䂐�@z�܌���K#����"O0��"��(Ј�j0-º� T"Obh�r�.+�0C����,E�̹q"O�S���|ء�&�$=�}X "O��R�?��[a`��/:� �"O<�;� �=��4�q�_�&��"O�XǤT�t�\A9E�ǒy�혰"O���N� /�0IA%G�u�Yv"O*c�&�t���r�B�T	� �"Oe��!�$9t��f�_�"�|���"OR`rv#LHH�I�i�4B�pLQu"Oڽ���� ^��E	�~�p��"O��AG
�>�>d��g��� �"OB����[�P��d� fU �=�"ONI,,��"Q�**a�*[�!�d�7:�d�V�Q�~�6����T�D�!�Z�A�ܵ��m�	E�bO��!�d��l2��#+�2 :�`��� �!���46(���J&P�y����	W�!��P�o�vMZ�B�|��1���!�C>^�X���{��=��얖o�!�ă�<ۼ�2f���I0=�JD�e!���(A�^� 2�Z�F�l�K��A��!��;wA�\�ש,H�� b�@5!�ϓ(����m�09�P`˽q!�D@�Gl���]�O��`g�1m�!���r5a%+°L{��1�Ơz�!�D
�;@X���N,�[���Q!�$O��$����b�ڠGX�,a!�f� ��X�~_�mA&@�$!�D���l5�#�JW���q���>!��/zV��I��mSԂլ��u!��^�rh����=q��sDMZ�Z�!��5Rz"@�����6DJ�Z
&�!�Ԅ8j  �d'�4D���F�!�$];��!4M�p���Sc�V$G�!����5A&O�R)>=q0$�!�d�6tF�cB�;r�Yc��j!�� �$c D�u�ʌ@�R�5/f�s"ObP�����C"��:P���*�0�`�"O�9�J��:�H�;��&U�
5�P"O���^XI�����9��"O��X&�֕F]�Dm��`=�"O�ŲEK�6=a~ɲ���!J�{�"O4\ɒ��-+V!��%g�#"O�%c�Òr di�Hج<|��"O�� �鄌uܘ�'��O�|�"O�t�/�R<p8���9�@��"O��QV�D�*>�h���"����"O�|Cq
�1�t��$i	(P�zM�2"O��Ы��)�q�Gǉ�SbF��"OB���  �   ]   Ĵ���	��Z�Zv)Ċ;R��(3��H�ݴ���qe�H~-�8L,<���i�n�?
.Q�0�đmz(�Ӥ�._6��)�4<�>��' ��0O��@6�ʖ���:"m�&To�pS�Y2j��RߴZBqOR����D^*�MW�[	A�Ʃ+oY�Y��,���V���D 8Qf}I�4$���.�응e�:ל�;R}��c��e�Hu�Ҏ��K$ ����6)<��'���v�Z&(%�OR�2d��v�4�
��ȜJ���ʡ��g��o�$�?i�'Ed���=Q�)-O,��U'J�D��\c�(y�S菳tT,hĭG�WĂ)�O>��M8�zrF�O�mےl�&�,a�fg� M-BA<O��������OH�h2CS"g(�\�-�A��$�r�p�'��IExbkN}�)�?-|���!�T'.��Q�L���W��3F�D� )�����%ߖSjՙ��ʈ.
��J�A�'|ZuDxR���3�|PS�C�����tf6yӨm�}rBK�'�N4䧭<�rME�{�X`�b�,v~�l(O��9��D�<��'}l8�Q�20*i���5g� \A"�V~�'�%Ex��Vߟ�	wA̙D���1!.��8n��X!.&�I�8��x��x����w4����4zxӤ�\.�~R��x�'��(Eyr.ԱtCDI�s�M'�`R���?i$�d}B�8����t��u7:���*eB��t� GOR(�P�H�ƇN�7D,�O�%���\�'}����C]~��t#��� g͌�	4��M>�d�ۈ*6�Q�<�I�)�Xa�(Y�=lT�fЯ�PX��'Nl��@ ���0 ]����91@r�1:�.�PBkӪdn��M��/>
(�%��r� ѹ�蚓��:C�i�ф��$ag*�[��ib0�!��#bЉ�$��.q�<l���'�O6�X�f8��A�dU���9���O����؟�y`N*�Mc���?�aO�� _�]�Ā+pu
$ӤW��?��F^`�b���?9�OF�n�7G�&� d�Dv}�ǒ�����^�nO8m%G%�0<Y��z�0œ�b� Ȱ��XE�'�_�l�v���+����=�����O��m����/��F��V�2v�t��͟l�In�S�O<�hT��|�P�넪Ӣ�m��3�rn��AK���g�V�s�F��?���	�����2G%X���eϹJ0X3���=W�C�I�Hkd��.&3���!!F�P   Y
  �  "  �  *(  �0  37  w=  �C  J  QP  �V  �\  3c  si  �o  �u  :|  *�   `� u�	����Zv)C�'ll\�0BKz+�⟈i�郠+��W<b�"	;YV�EnڕGM(��T�GU��*e��1�f��A�!s�#�uE��ݹh�ʐ�ӊA�& ��L�̀Zm���z�ƛ�(��s���C"`���埳[{6�!�D�.�H�k^w���Y��O���d�� ��6.�t�Ջ+0 �0P�Bi4��ē��mM�T�O�|z��lz=�W�'�r�'�R�'�P�2u ie]P�ka�B�Y&�'<B�'�N��!_���	�E������
��&��'B�Y���R�5��q��� �'�'��/V��Mk�'�-�,Np�xgI��sl���ѮN�uўD��>L[�T���:f���"[-��듶y��1	,���H��v	�v��I�E�JqKr}�� �O>���O��$�O�˓�?y*���]Od�5P��1/6���?q�&�dQ��9�޴m ��	|ӌ�D���Y�޴,!�VO}ӆ���3h�ܻi:2���Q6!�:)ov�=���0r���D�z�� �W)V�wܒ �Wa/F�lAgHU0u�ҀnZ �M�i$��՟�i��ۄm̔TR��!���� ^9/�d�3׼i��]+d�9t� �g S�sn�E��ؽ@�Zc�!`�<en�!�M�w C,����HT8'�p���@jAr`	o,8��\9��6�a��l���mrT���S�d,yp�H81
�( ؍�C�S�GvF}`7%إ#���"��286:5qܴ{���hӬE9�nK�!�<p�;D��I�E�(M�T���bU, ) Љ��
�܌n��u�Tl��n>:���i!*�	Q4`	��^�� ڀ�	�1N�ёJ�.y�e�����'���'��=قuӶ�d�OXyR�"��?+��"֊Ɔ|�h�@���O����9D�p�$�O��S[�f>�aa�P����`��]�4�����E{�=O�h#ܴ.(���1�/��$���b�Y��F���6���@�axRc�
�?Q���DB=t>��r����0�� � ��'�b���Q��� �\#�<�	b���h�^���#�l�8r�� �+Գh5���q��O�D���&�'�y%F	������ ��V�Ԝ�y��2�d()�C���)��2�y� X�N��H���z����s� �y�A�LdFz�d@^ �s��y��=�j�@��7�����+
�y��(�q��*5)��+#�
�?yՀ�~���������(���J�f����$�(D��oئ18(�B��`%Y�D'D���f/i
�c`H֨b�0a� D�h��Խt��za��<q~��F$D���W*E���a5��MӚ��׌6D� �C	C��}�F��f�a�ɿ<q��g8�$g�������%%gI.9�H1D���$%��y*�H�e��3�*�X�C*D�D�RB�G�ݛÃ�0��� p	(D����G�0,���)A�d����%&D���D�6��w&�; �n�hϓھ�����V&3�4���d�!sYb�2%e� #ax����L�jM09�(���]��|f��|%�|�U!�"پd�����@YT-Ey�@	EQ�0F畺2�r��L#s+�cdlE>\��D�	���A����8g���Dy��H��?�d�i!l7��O�yRꌻ�
xH�Bэ4*�8ѫ�O����O|�d�ON��:c�PsP����>�*S��|Z�e�$1�O��	,8N��p��%'�L������d;�	¦z�(6��O��ݨ'|qa2aB�g4 7a-{B�I�k+�,�@[�.��]�'�Y#�B�I�Ul
	�g���ʐ	BD�V4�C�	/K%��ф�O�2(�2�;R��C䉶�]/�Jl�#�C�4���"O:̉#��k����.Ĵ8ՠe!��c�l��On�dͳ�th$��O���O����b�h%��K�9���l>U��a�FJ���""@ɦ���f�?_�zP�Oo��xsdΗ$�bU0u���)+ Ź��?v���sB�z���A$��+2�c>c�d��h��Ե7o��3n�܉ ��O�@�'�ʸ��bY����'��tg7o�nY�>}�x�@֯��"O: @Wf#'�~Y�bN��\���X�� �4���|�O��$\�E�!L�z��	��T�ht+2�I")�:�)��W����d�I�?���쟈�'�ҡ�aL7Y �`�G J0=����&��Ȣ�@?Ohp���kмZ����pc[H�I��[
Ɯ�N�����	�z!��q�����4�ME��L4��4L$ɔ��'oS8iB�yp0�'����~�'`�Pp��-�x�i�*x�
�'j�hV��.?�*�p�咹f��H�I>�u�i�BR�d�i�,��i�O���ANNjٜ�	��?!(���#G�O��DO�L�$�Ot�S�]��<��&1ePe� �Jҟ� ^�S��4�r�9 �"�����'p�u fm��/9P�醂;��_�4���P����Y��ӳ�0<��OD��H�If~�љhrl���@9�j8�����0>��M�U�X�`���@���p��a���a��`b`����19���	�JPN ��Ixy��/F?r�'��_>5�m������)�+>L>�r1��*m �dȟ8�	,?���s�Vk���L��
�ߟ4�'9���[�+��`G=}t:<Ir�=?Y2��M���I��ˢ	�Eb��
:��r���)�<����e�!ZdLûb'�"ѝ��[���O*��=�'�y��s��}Z��M�^Tb�P� �yb���<��8�$�Z<,�L<B�'�:��OiD�t��/WzH�!d�K��A���I6�V�'R�'n��grT��'[��'���^�|�BC��=1����_�1OTY�R�''"�#�J:|���i�%���f z�y�����0=q�����w�q7��i��[̓r3����T��Sɛ�Js�2��Pl�zsG$D����T��e{�I��+D�h�	��HO�I/��ZT�}�G��jc���"ڿ'S�A{` L  G<���O����O�y�;�?�����$IO�_�f��	�L��x�jF�f�hw�J-� -��L�� ��yRn��,��T�&�!z�s��M�~2�IÙ 
R�����0=��ጔ����Ej�Jd�կ��N>���ٟT%����۟�?1�a��8���I�l�;|N ���С�y���&R\�usU��VW$I���X��)����'A剴;�DI�O ���P�"D�Q�@�k혠�ʆS=��$�O"����Ov��`>U�"��t�\|%�� ƤULH
	9I�3jS�5�q�:O
�{!�D�H�r�O�uqۙV�DBC�ւ-���SB�'�̴���?���?WKɐG��T��^%�m �b����OZ㟢|���9+�i��H0{��M;�l�R���B�{�(�Xd�G�lC<(�g- JX���PyR#Ũ9��ꓵ?)/�@!3�
�O|�b�唘.�4qKW�ߐQ�r�"�n�O��Dѣ@��d�7[�g#U���'����8E���h�C�
վ}�a�_8S��I,!IN���&��I�5s4.]B�O� )� �BQ��Kg���
g�[~ŏ��?!��?9������ׅA�]��E`�T��\��&�|��'�azr]A�f�
P]�R�f�Z��V9��O�\Dz�ك	�hq���Ly8�2gA
�F%beɘvJ�O�剟\
�`�r�އy���۲��"H#D�@�P�
Ax(xq��K)��9p�+D� A7���!_j�j��M����-D�ē�
Du����V$`E�A�B*D�X��*[�O��Paψ�m=�*��#D��nT�o�fT��,�a��1˓�<a��M8�*��!Gb���ǒPh؁ f D�@7�[�L`p0aQJl��[E�=D�8#��O'U���p�\�8dTQ�4�1D�\I�MU�A{�Ԓ7�M6(��%yDf3D���%&還�ю�0
5+�#�O����O�5��Q�&�V��E�5ZgRA��"O�����*ID�Q#�	�\?�<�g"O���H�)i���7��r.�ЃF"O��ӣď�{�5m:���P"Oph�u,���8��Pc[�%��"O�	`!��@Y��3�a�)zr����I���~�r�D�b.^�c�ŋ
D<�y��k�<��	���{��y�!��f�<��ԌV�e�Rk�?x1Ne	 ,a�<ɀ�Ɩ)�aK�I�����p�f^b�<�Ǡ"l�`�ʠD�1Iq�L���H�<�4��;8�r٨�IQ�z� �c�KO��@x��(�S�O�d9���#��%��X��B"O�lk�J�CʒLb�oW<`���BT"O2ȣ�S�Ba��-8:T:d"O ,�!��}�����uS�"O�#�*lE�x��ڇ���!"O����ē	n��a$�J�<�2l��_�D*�i.�Oj�Ɂ��|��8q6"R2?vdJ "O� ��Y�.k~!9�̙wQ�
�"O�mr����3)TŨV@��#�"M�"O]���) Jh�H4/�}�<��"OH=�
[�dCRx��W�-p�s��'�f���'�>x��ۊN�F���N-��a	�'��9�E�b_^� �C݀Wݸ`��'C�E�ɌDv80��GU&@�L���'o��X�����$��nO�C��հ�'$��R)�Y�� ���(7�f�{�'�h�pd/��t����7�Ѹ(-�X3��$��e�Q?��E
+>���kn)<�rk��$D�|�dL�6����E�P�,8�`-D����˞%	B�3��O�3��0٠�6D�����cPDIqa��W���6D�<0�Dba֋I�7�x�����Ox�B�I�jS�8�l��L�N�j��ܕXg��d�?l6�"~��]�O^~9��1PNM0�	֞�yR��3p���Q�� �L:fA2� �y������)��VC)���'>�yRc_8|����*@��e�&���y�آYb��UL,!���2u�A�yҁ�C(���P�"��CWcŊ��$����|JC�B٪�hϦ��̂G��0��[�N2�
ݰZp�4�Z7G@��������MV�_^���2o��.8�݆ȓ$��1�֓;�t����/��m��.�`Q)c�ںfv������mvn�������ɻ���G�J�$��<Xv�VRB��9>�И���M�x�ִ� �
.]�C�	�ZM�4±IY;-7\I	����g>�C�	�>�č A�ŢW���"��,��C�ɦZq���D���{���`%�	�x C��!M�n��BkNt��])�%C:}��=����K�O�t
� f,hB�,q�����'���YR� )�<��a�n���'������	��@8q�T<^� �K�'^:�+�ʄ3�D�Q %�e�~��	�'��P�d��.S_V��J��T�~=��'��Q�G���i���GԂ=�>���Ex��iлI�� 7�9��E�R-�B�ɍ>�֜
G��y+H�JEA�SnJC䉱a�������.�7�L*iZC�Ie�`���ٚE/J�X4	 c{�B�ɇ��`�6�X7Iޭ�$J-I�B�I�P®��p��gqƵ!gH��k5<˓G`8��	�n��uⳎ�0���ӃB�Ob,C䉰-` %
D䐙h�4�Ѕ��*C�uP�p�4��%r�Z9"���w�B�	67�����j�l�*���T�LG�B�	.XfU#'C�5^ì�ʦᑤL ���N3��D��n��D�B�	p���	<o�!�d�2'��P��SBT �P#P� �!�Ѥpo��K��^�(���7�!򤒗�8�z��S+8��X����!�ή#�����@�9zz�4)1)�j�!�#e焸Ǭ�8i�h�3e$wў �4�&�'��S�ݳr��xy��k�����*��5���( ��M
4k��ɇ�Q�>���]|.�	ñ.�0U����(���`%���AAF�(A�ȓ'�:�"����s,6�X�}Js"O�$���16��X�lءs��}���'Tᘌ��ӻ
F 0 �Ö�J��R,�p��&���;�A�Gf,��
ԾV��X��S�? ƴ���?5��\���,��u�p"O$��W��Mh�JL��:�J<K�"O� �� ����P7k�,�h��"Oy#¢��g��ؓs�A�(Ղ�ےR��ɔ�1�OΤ�f��� ��Gʎ��"O���ՇʶC,p!�z̋T*O ӡ�U�	�P�G��VT(�	�'0�	s�`��5c�tIG��:��Y��'�<��!��/I
X�F`�!,tn]B�S�����a@�@�*�"a��1�V-��8۸$�B�\,�#)��"	�9�ȓ<|	s�c�4_����N���ȓT���C�� 9O0U�!I�)"��i�ȓ	�� $	�X���M�(����F����Û�Uܘ�6 ��؅G{�a�֨�������q�l�a(��&p�"Od�`��ro4� @�E�pm�ِ"Opa��9��%8B)?|UB�"O6�ӌ����ū�-�i7���#"O���g�I6BvD`L؞m}����"O�9�hfP!�vAGu�1�'p������#mOF�ȣ�I�J��(hR盜/h�����iV �:I{b�2;��B��;(���k�u��`[ 3
��B�I�9Cf\Z k�=s���e靰-fB�	��r�{��[PNȹ���I`VB��7nS务��'��8��n�'�Lʓ4`����# U��Ń�';	+Ԃ׎_�"B�	3&�`�3�߄m���j��(�@C�I�(;�;���.!Iƴ���ߏ9��C�I�Kj@��	B�[�^��n����C�
�r���O%l�y�#W�c1���Ĉ8����;M$���-,TĶ���ы�!� ��r|1�O^�kV2��v��Y�!���3^�v��ѥL*!�� c���!�DĈ"�<m�#�Ƶ8�$<z��Q�~T!�dZ���9��n�V�\,s"��qr!�
�� Ց�e����@�pK;E�ўP��:�C�V�����P(�en+�@C�	=1gH ���7k��ЪW#Hu�C�	�'�L1ॆ�_���Q$d�w��C�Ʌ1�����Ή@���rDI"R�C䉾qT��q0�@�vl�`[���3�HC�I��)1wIW�Q.��7��^��dD�h�"~�(N?KÒ`�rÐt
��R쓘�ynoԾ9�&�H�7<4 �Ż�y�e׿#"80��m�2���Ufф�y"D]O!,(���X8Nb���̐��yB�<9����I�f��d$R+�y�(ȮS�:)q�B�\�Jh;$����$�>o�|�!�NK���a�C���a��V��y�+Z� �i0iX�h�|��"!��y",�êUۂF�1d�r�9�y���d���0����a�)�(�y���Fk��a ��
��#CΣ��>1Ԭ\?��ȐV�$)��GI�X͜�I�J�<�6� �Đ���.&���JE�<	W �*vw���.�}�\d��eH�<��I�q�v�FJF�$�V��e�C�<Y1���j�5��O�V^¥��|�<	5d�f,\ #�\��x�!g\B�'����iCJ
���a��&\��I+A.2�!�dA�BT�����2xp=�����!�dD-J1�q�ͻsl*Z��=�!�� �Tk���'%%e ��y뤝�"O^4�V-�$�pQH�$�N͘4XT"O�LX�!���=��@Y/b^���'�|�����yR5����8�E��N+ I��X2&�C���}F�R�}d>`�ȓ��=A���B��� ��S!h��ȓ8Ѡ�:�[4w $��ߨ#�Ԩ�'-�qG,=:9d� ��E!"6�uS�'�~���l'?�v�Ka䅼b��+OA ��'�ʕ��$� ��q�3=��1�'9�A�#	�Ve�%��\�m�%��'��<A%ܠb����c�q`���'����I���Ɯ�D�@;z�'RT��cI�<��u!�I��p"> ������j��7"@=��)���/�̅ȓ8z�[�C^�s2ڽy��6Z`���p�g��TN�A+�d_.��g��'%�>�Rŉk�hM��
�^�H�!�7k'F�j�BG�$()��o������!�dR������E{2��˨� ��)�!��@y���;��"O�S�)>������ST��Y�"O�]�'�՚hl$U!G���,���A"O�L���i�tȂ��\�_ò�*"O, Jŧ�O�`,���Q�TLJQh�"O�h��	2H�D�8JL�H4r3�'�b�x���S�!��щ�e�5 B2��G�����>�rW�;Z{� ��2�v0��.���&��%b�v&݇E�.E�ȓ,��HqF�B�P����]JN�E�ȓD��1���HȖ}�Gڻkj���Ɠ1P�[��8����(Q1 �@hȋ{��ؐ��$F<vy��'�ҙO9�TB�#� vfbm{�M�
$.�8��^&\����?A��"i0����I "Y�2k�>ͧY��T �HȅU�y������D|2N]>Oĉ��X�>���t����T��š�C� [\Q�2��/R����Ob>�� $�p֎���.��gD�<	���=)Ć@l����.��5�����I��)Ĳx����{�����R��9��Iޟh��O��R%e�
	簥b��Ф2GDy�3O61���16���Ba��o}��I�#�.�۳�]�J��C�L��"<������.M�2�,է��Nu%��<	f�P�gʁ(���0�;O ����'Or����f�~�	X�j�xe��Y!��$T�ȓ���Pc�nݪ��鉴!��eF{b�9�'u�"l�����N�j�'�]��Բ���?a��E�^J"O�-�?����?������)48{PO��c�|swL@�������Ω0�TՉ���V&.����̟f��>IAr���҈D�#&��d��'�ٗD�(�6`�$õ+O�8`�?ѱ�4�M�R�������L�:�)Sc1)���K��*?ic��֟���Y�'d�½h���s�T�qF2��¢��mD!���!X���פX0Ѻ�ȑa�=�"��|b����D���r	�@��&%�#H�"6��y� �OC(�	ҟP�	؟���Ɵ`�	�|��W�v�RԙvmQ��Q�Ūs޺	��Z�&V܇f���B�	s��h�4K� q&́z�)�n\Tr����D�fP�A���6ǅ>�Mش��O�H�'������3S����X�f�"��'�ў�F|r�J�}�t�$ ��v��k���y�΄�t�z��AoI"E>i�fD�'���¦-��pyb�5��'�?�O@`�X��8X�|�٤�ٔZ�:����ob�����?���t�D���0i�<���e��]��Ou�5�'�ٰ�fM�$ y��ȉ�Ą�?��g$Ф-��4�é�|�� ^MJiq[��:��I)w�h">�4�����	Q̧��y��Z*Bm����9����'z��'A��h��#X���z"�թHlJ���7��C����^ s�V��g�M*���q��YK��io��'���78J��	ퟠ
���=��9�q-H�)q�	�'�㟘CïԹ-�������gb�3�S���\#T�t��c��9:����F.��$�,6W���rfO ~ٴ �"0��W���F�����Ǒ��� ͓]�`������'��� ��P���-��d� ��pW����"O� 8�%�9���"��Z(@3Q�"�ȟ�(���#@v��#M���vQK��O���O��A&�I�=����Oj�$�OrU���?���6v�	�"�W?d&v��aN]�D�d�'Q�=:��J�*��� ˟�h���4�8Z�柸9����>h`��I7t 9��\9�@�g�'�h��C��[Br��`��u=B��O��*��'�b�'��O&�S �u���L/ (ЛU�t�,B�Xdh��aŵTfNqc� A� �2�d	S�����'��	�2$���AcH �ࠌ>3C��F�
_4��I�����x�SٟD�I�|B���-f�P-x�B��%p��'Je��(�'	�t���ՙxڷ�I�=*)�	ȯ	�$L�YE��Ǭ�0sִ��<I2F�P䉞3�M;ݴ��O@�kp�'E�IH"�_�V�����m*`½�G�'ў@D|R ��X8� �&`s�됡���yB�`�Q/b&�"���S��'2\7m�O ʓy~��ܘOI� dK�p�,�a��}����DC8*sh�QV�Ԛ6���S�K�!X��0�(����En���F�p�o�BG>9S�򄙩�r"I�+��q�k�{ ��R�KZ*+�J\�C.N�l���,�AGz���1��'���'D�鏻i�8;Ug�2���Bbi�l=��'A��'��R>�ExR)�af��q& .��S��+��>Y�]�x��k�GwnD���2-7�K�
�<���ߛ6�'�1��X�`��hQ ݹ�dT�ɾ�	T��~�	T�'��,p�	̵3/2Mz0L�5nr����iU�'�&5�|��	��j�������<Zv ��CHG~b����7}*��$C�N�T쫃�F�9i(�9c��;EL�q�!?�s�>!���Y�$�x�Ӵ&���"!�(פu0��
2|�]cR�>�p�O�}�4�B�2 �/1��<Zf���i?�ʕ	Do�dTq��K� A�t�S�e�@����7Sș�a��'�������wCEE�"Y��Vi��y��-`��1$e�oԆ��I9��I)V9�'�z7풳�~	�悗P�d����X�I�_��'�,#��hG���qb�Ù;�&1��ϑ;b�dM��S��'d����O �R'E�g7��ZA�=���;�c��uR`� �@��'�j���'C1��i���!�r��$�F�|����q�'����8����9O�y���O q@1�P�W
��3&AϠx�(�*��'Vi���/z�Ny �G�i=6XwCH^��C�ɝ��=
%�ްOt,h��j��&��7��O2�O�1�����|n�Q�leY6�5,�x�g�JT:��䓺hO��r��r�)��=q�턅t�.C䉀��h	Q��<v��i;0oğpC�	-uɘk3(�)+9���u!AK��B�ɿp�*E��-,_dȋcg���B�/G2F!A������@O�d�&B�	-l�,#��ޱH��i���ʬK,C���)��%�Ir��D�ȯXK C�I�=���«ٮB3|U����=�:C�	:�$�����U�X)Q��<�HC�Bxe�$t������ؒ�2C�	�_l�I�g��-�p��\>�C�I��S��ۿ�c�-�_�C��=`ޮ�+Q��z�6�)6������2��аxǬy��" k�:)c�()�4}k�M�2f�)���n�`�)*X(|)�Ý8x��ƈĘ(�Z5���?JE�,h@��Z��<�-W6@ȉC���Ik�a�!�Of� �h�&]jT�u��+z�0�	��u!�)f4R����7(�lQJ>���$i2���B��bO�R�FC��>��p�BoD�(�B�;&��?~ C�	3ˆ�@�yj"5��"�\C�B�I�?wش�+˯i�	��G��$��B�I1e�,Yp��R�4��C��,2ZB��6^�
x+a Y8@�`'��<�,B�	*.��x��鎑PH.��g�B�
XC�I�!ZJ�hsIA�&��KxC�	�B�ڠ��<��e8kH��jC�v��9sҍN̊u�s��	j\~C�ɦMC����+�8��E�[�HC䉿e�4��q$B/4zIt�D�@C䉻JD�+�*ϪQc�xt�ߎl?0C�)� |�j7�\.�qU#�'� %� "OB� AB9�y����jM��"OpAe�/	�y(ACN*N=��R"O\��w��]NЉGA�Y P�z�"O�D�4%O�A�ZP���N	<�PW"O�iJ�G@�FnT԰���3V<�P"O�,�b��h�T=���?"�����"O��b��8�.�bc߳8W`�g"O��ǭ(ղe0��ۈ ����6"OLA�7d�&m~�QBM�V�R=G"O&8��,R���I.
�5��"O����L�%�|x�6'��f��<�5"O�T��ހ|�����Ky�ĉ�"Ol���ȓY�L����S�.�4�"OvA�T�g�PcIݸa� B�"O~�I� �0Lz�ȵ╭KЌDu"O�hwe�b���2�x��f"OR�&Ѩ-2V� �ȥ1�ti�a"OT��V�06���!��.L���"O��{��ѠDri``��:�d\	�"OB���%:$�\y`֏��f����"O�l��M§�B@�T ��#��L'"OT���5%V�rPn��Y}6�X�"O��bzI*��(u����e"O
mArF�+<��Bb�#oh��"O>�q��Xy�����I	uh(r"O��@�����JH�^x�!u"O� s��5"���C,P)��#�"Oֹr�ʗ�Q����� �B�&<+"O4�1��sL�31` �Z:v1�r"O00;5(ޕ���@�/;4�0�0"O�|!�又}�<`��$��.�t���"O��p'յQtɠv�GK��li�"O��el��m��MЃ��+�|��3"O2���A�|v&X�B��My�iW"O��a��=�Z������<вp"On���@1����ք�V���"Ov�;�˕2ςM�1��`�(�A�"O´qB$)%��A���Y�	 �`@D"O�9)u�_������@8ؔ��"Ov��"K	�8q�U��u/��C�"O�ш�,��E��Al�v�$�"O(����A�_}L��k1�4��"Oũt� !ɪ���_%���8�"OD0��5A�P�㊏<}���"O��2��$�6�H� vF ��"O@��T���趭�5t,�i$"O���e��UK�Z�iW�u��"O�8sL�	:1��?>,u�"O��Pt��-X<UR񲢺���@�L�<1R��jH���P��,�j$��&�s�<���QIr�HO�@Ǟh�Q�Z�<q%!�8F@\����nnRd�GL^o�<� HC����D$ϻ�"��B�<�QB�V1�lӒj�1C���:��S�<�E��]ꐜ2t�G�s2�P�<�2��m��e��@�5y��r�DE�<�oD�# �}�R� ({ ����<�E�V���	'�\#�Lw�<	�)Ε]�8�@�C��L_�#��t�<١��f���"!�!u�U��X�<��ʑ��u���s�z�TM�<�E <�L���̏R����I�<1��[8�B�2�/R�PI H^�<� �a�G_�hB�E�5�X�sT�|Y�"O��C�jL�G����&-G4Z�"O|�p�O\��,���>/T��"ON4��J�>j��HC$�)`�!�"O�a)AG>D�zw�L�u�"I�"O\y����E�2i�i�0�=�"O\�9�P<��v�L�=�@�"Oֵ�e��1	I|��B`��C�m �"O�hJe��*�!��͋�e%�B�"O��C�*B�[��1��~��:`"O��B�6��Ċc�ܰ\�,� "O��K]x9�J$�$|�4�"T"O���$�6�|pH��+����6"O�I���'��)�b���up,��"O�葶
��i�Z� �̞�6c��"O��HǍGC�b�У(��Je"O�ts3$�G��rʒy���"O�0�#��(nԩT�1'��(S$"O�9�:sQ� '��$ ,m�"O�ỷ��h8ii���Yڣ"O`�D��$c�(];��KB��"O|��@�d�֩[������u"OD�ذ��j��k-v舰X2"O,�곫A��M�P ˊԘ%	�"O\�jC��_:��s��Ǧ�r|�`"OD���-�E���.�_�5Y"O�M�T����,9��@�b�5�P"O��H��!,6��Cl��c�� �"O���"'�9k*�X���ؐ��EQ"O���HM��0����Y���P�"O���b�����7@��y�C"O�4��l��8P1/�'ⅉ�"OB��TDۊF�8��`����H�"O��s��ja�Q
Y �>H�!"O�����zמeI�nZ�?���SV"O�\����!HX�pCm�F���"O�).Ӟy4�k�.Rؑ�"OJ1�aZ�nx��쁮,��(;�"O�r6�� gJp�;�LB�r�sC"O>����ڰ=�2i@"���~�S"O6$����2���`��C�9��h��"O��C�
L:a�&�R�Eڕ`�����"O�X��F�)IMN0Z4F��"��D� "O	BoR�cA<�E�V{��q"O��A��Vs���ذfD4���"O`�	�??����"C�*h�!"O&�1�<m�<���BA�t�:�pU"O�J^-@��v^-G攀т"Oa�d�D�
��$'� x��"O8�A�lUf�h9d 8xЌ��"O�Q��O�C��P�sݤpQ�"OR�H���h$�5��cڙG�}��"O�+�녤c�n�pç�+z�*qaT"Op�A�CѺQ�"aK���F�j�3"O����$t�^�0�e�,u��=*�"OFL�F��3cs�!�g/��8h~�H�"O����%̮L !qN tp��E"O�S����@���`�\�S��ī"O���ú�a�qnO��=��"O,X��1Z����&�sܬӆ"O9 0JP:$�Ԩ����$gR���"O<A�q�Pv$ �U�F��[#"O��)1ϗ�4���(DA�B�Q`"Ot�(���z�e��ز^(��"O� ��`�q�<�s�R1%�2X9�"Oii��4=rE�0M� 9jN	��"O�ز"D��e��hu�Hqc���"O�<ȁ�T�]��FkW�\EJY#�"O�A �B�'�D��S>-1�H�'"O�Y�C�x������*�;�"O�遊��8YX�`�F�n
QBF"Oܘ�5��F�
a��$�FYpt�e"O�=��㊸+���3��{O!c"Or(AL	�A+D k��R�2��8�"O�I� 	Nt�h�š�b4(�"O�,��dΆG_�EZ#-��P���Z�"O$\�$(ۨph����"�!(��c�"O�4���J��Q����a�~Q��"O�1�(�!S��B�o��xl��ʂ"O�z��Ԅ��G��-&���"O�,��#u�Z C��';�q�S"OB���!�ՙӄL�6!^��"O���vmI�3�	�uJ�be"O�C�$���l��G��3�\�Y�"O�t�%/��r�@S�d�>z�D��"O:�#@�Ѝ�&���2e^�"O2�`F@�+\xe�&�ԕ%D��"O
|�`�a(�]��Ę7Y���"OZ0a� �;jX�\J���](@���"O��sr� *�I�$萗\#|i�"O���Kʹ%J���ˤHj|�@p"O�iٶ��|J �����N�̊�"O�=��6_�@�*���U���h"OҘ���H�Ig�(�!�*n��8 "Ot�HT,��G�R�`�T���36"OHE
CkB��HB��*"��"OLQCʃ$6팀�"�L�!�aK3"O Ց�N�E5Ԣ&L̂*�F�@�"O�çI�jI��1�TV���(s"O�4�%���g0����
/�>��"O�%Ǒ���|��N%��� �"O�XP%BI�b�^)��ŀ�i�,��r"O�ĸ�-��E�"��vjگ%6��"OH���ͯ�: 
�� ɜ0�H5D�tp��Ud�x'�]�zJ`H�4D����!:�R]9� m0�`�?D���/�Q�����ߌ�X�d�)D��*1�ݣN�D0rG�!M<Y�G)D�@h�)��C=L�z��;eh����(D�h�d�1h�]�0MX2"���A2D�l`��
5l>,B0�H����p 0D� �u
�d�RC�gF�z�����-D�,K�I�&��8�3�
I�`��*D�`�	��<���6���~&��A�;D��
¤�66�P������腐0�>D���"K��5'�E�A˝_�!��>D�4�$�ψf�DC���v��QRV�9D��#%��5���� �>e��P��:D�<X��\g��8[��B(��""=D�H{��K���b�_�K,�4y��9D�p�%GŕPp�hФ��2��H�@�:�I�^�T!V��>j.��QB�6%ր�O�͹�$U�3���T.=~���"O�d+�A�}�0$�D�#Ef4!�"O|Q{qm	7F�Ĩ�S�ʪ
E ]��"O�E��9���H���"O(1�2ˇl���r㓹va�� "O�}��"�s�����_3�Ѐw"O����� vS�m�p�H�@(3�"O� �D���C�6���A�6�-��"O>��2�F�#�[Saj�9J �X1""O<ځ
P����؁�³<߼U��"O��#׎�&Pg ��Ҁ���@"O����صRZ�a�T�L&vܠ�� "OFu�ҎÚ{#:%���Qlڄ��"O*��2c�)\�p+F�	�2t���"O0j5�':�؄Dh�e�V8�y",ٞWVrX��%A�H�๴n���y�Ș�aF3AO�y �4 ��J!�yR�C�T[@ej�.�oz�:��E��yr�W�U.(�� �;j9�pq���y�$�9A6&���C�T;������y��9��XK6g�/F�f�v�;�yd��\&U�O�4��i�o
�yR�K7],�ЁE�A�ym4�s#i���yr䚟&L25Xp��5uF�� �¬�y"�V��^�r�GDE�����&���y�O9�$m9楁=vO�A�D%֢�ybK��Qz%�V�v��1��I��y��φ+B�m�'��m�v�2����yB���_�f=�AjQ�h����nɧ�y�$� vP��1.ń8t�l2 ����y�`���ZhԀQ���aڀ���y"I�)j\b����a0W��`�C��"n,�A
gH*P�j8 1Ι�0�B�	:9( � �^77:@�r�.�B�IN�1Ѷ�.t%,��5S�d�B�	!H�� :���;T�X=�%��57��B�	QV(|�B�
nKrܑ0�[�<�B�I�:VV�� Ub���';8���m�j���`�.^�3`�`	�'����`F�a���c�_��d��'�,Ȱ��~"��׏�=�M1�'^8u{5m�#�9����L�l5q�'Vd�QłD�0��5DE*7(��
�'aTM��!A^~R�U�9�*��'���kq�N)�F�z���&%��"O�d�Cm��mV�����
c&f$HV"O����!}~0�çGK�c|0Hq"O$�e��2���9����N��Z�"O�y�W�A�����
�!�~��c"O4q��Lqo��#�i�jg�}��"O~�ط��;����T���S�ΜJ�"O>H�e��',I����V����"O͉���gh܅���$�gf8B�I�'sL0�!*�tQ���U��PC�IA���  ��J����O���B��.vu� h1U� ��.N�=�C䉹/��� ӯ_,4��%)!���C�#,��(�.��1Ȥh4�L3�C�	6;��I� ͯR����Q��.wjC��){��@��9-b)3̐7!*C��

E�X��b�5�����o݁uԴC�I�Pub�.HwM|�����C�I�
�\��� �x[<@h4�ҿE0�C��&w&|�Ă�4;4�"�(�RC䉉L	FH���U����R�^��C�I�%�v@s�	U�=Μ���:l�dB�I4��)b`���N����ɪ`��C�I�PB�A�kH��:A�A㖯P=FB�-#@�
u�IM$����;p<B�	�VNdP�t�	$t�.]* n�=B��|���h��P�TPJ��	�� B�)� ��9r�64ȸa{f��%Hċ�"O�M��-Ԋ:��lyp!ۺU�b�K "O�b�E�m��9���2ϖ���"O���ȺsZt���ͽ,de��"O>��AIM%��#SN�y��x�D"O�`�u�U¤�2�BB/wN����"O$�b@�<%'`5�w˿%����"OЌ�N�4 �.�R�M�/?,���"Ol &�L�Cz�jvm�Dc���"OJ�+���z�f ��4P�1��"O���P�s����3b�2��с"O$
�a��P���@���P��q"O(T�E���)�� �*U��Q�"O�9i�<��(����!�beB�"O�	6�/xm�c��+:��8"O����Q�nn��0%I>�JAps"O�lڣIׇFI�e8@�Z.��u��"O��سŔL�X��PlI:f90�"O��2�׊
>0��',F�H*I��"O�օG-����� Ė3�:�Z""O���*ɧ9Kڐb3Ac2��"�"O>kVfT�_謄�"��Q$��{�"O*� %N�D�p��zx`�"O��0��.!M�%��=)�R;�"O�����ҀK�L))�"ќqa"O�8��hɅN�|p(q L�H�AP"O(r!�Z=Q˜dxէ�=^�Y��"O����	���5`]�6��g"Op��ʢ.��hA����
y�Q�"O
Ik`ϥ\K���V�wR��"O����S11�D  ɍ�4z�Q�2"O~����d�V�Q�����j"OҤ��L �h�ɣ�ꑸ4�FMh�'~Yq7�6������WZ��Y�'O84� ��$$z��[�_<T���2
�'!^�j2�����аu�҉��'�RQ@T-ܣ�W=oF�`�'U�(uc@�za��DȚk�r�H�'N�;cKiNfa����e;p��'��尐AAj$����H��c�'����Âܑ]�T0��U/^��A�'�h�M�,~���X��73��X
�'cι�ZhĢ�J+y�h�ȳ���yB
m����&��m�S���y�N;4��Z�h(&��(3��.�y����H���!�&]��g���y��P8��e�G��Jt΋;)�,C�ɺpk�p�A�!#�`���-�:GBC剳=�\s2�ȨI����+|�!�䝜ph�#��àX�P� �j�@�!��B����46�=*��Nx�!򄂦S/�����<!:5qC�z�+�'Pcw
��R�6�Sb�8L4���
�'�Zͳ�C�s��r��&`��	�'q~�	��^2g2�Y�+:�Ќ!
�'�x 7ުz�<��0 E�<�@�K�'�``i��[�#CMB�CĐ53�%��'�����KL{ �{T�V�4�"!��'Q���*	�]���*��2
�'4�icsFC0z�>%���84� ���'�T(`��<*$���A2V����	�'Ϫ��ā\+y�Fh�`��Thت�'�PZ��D;T�A� m����
�'��0s�˓�2�a�'I�![?>��
��� ���Av0���j�%�"OB貤��XߠQ�a�ށ�r-�""O.8��"NA�y(��w�tJ"O��! O>��u"V�DU�5P�"O��Y�8� ���p���"O�a3脬�0��7M�"D
�"Ov5��W�j�lQ�rA�^��q��"O�\9�i�8j@�:ǭ�Q�0��u"O�IH��53��0⣂���d�w"O졲�IǓ��s"L�9�hh�"OR5��Ě%hʄ��A!`��|*%"OZHL��l�r�����"OeU ��.@Lx;S�ג5>����"O�����u"����N����;�"O�IKS���i���j�
��u"O�,����r���1�d�455z�3"O��sB���X��8��E�s>�b�"O�UӒi��nE��"!`�>
��{�"O�0 ��*	[��s�'�4��!w"O搑�hD�{�z��Qmضz����"O,<�F��714��ЬP���H�"O�ٰϔ�\`䝳�c
�O�^iK"O�×��,mh⍳��Z>���A"O�c �L&}�Tc�Ŗ
�2D+"O�DKSC��T�`k!G�։��"O�	#/�:$z�̨��%be�i"'"O2@P�è<A���ui��"Od�lR�N<�ēF�ݎo@����"O�����H�������@"O�=���ר_3�
��
{�����"Ob�j��

N@䩐=a!�{	�'�#ʙ=iK�IS��ĥP��
�'��횠�

Z�Ep0X�N~Ix�'��$Pf^'9(���| (���'��Ô�"xtl�'W-m�Z}�	�'��1�`��C���a�1]b�	�'L0�(���*�4g�;/йH�'O�����\)ab�F��v<��'��,��H&,I���L�5�L��'�� ����
������+���`	�'x�Y%%աJ�������{�f� �'�P�zjÈ)�i�Wo؄t���h�'��<�HM��r����f�B�k�'���	���8HDh(�p�A.`���	�'P��ĉG�"Nh������'Dn|y�)�:���VJ�{ �'o\(1����2��U@Ճdz�K�'=���@ ����������V���']JM��@�r��9�*�	9���
�'� ;��G3B깪0J՜y�D��'^z�������~AA�G 82`R�'���Q��-@���s���>+��(�'AD�5��b@��g*)t���B�'�E`�霼M�u�&I.�`A:�'��ds�k��i5����B���$tR
�'�TyР�D�j�ȧϚ�!LY�'r\��#��D����G�?�\1	�'p���V�J���@�2P��	�'�P���?|�>�� G1Ib5��'K�y����&hI� x��>.�0�'<VM��eF�fY��* G�^BŚ�{�����M�n�=sB5ʰ�_��a���z%�LENݨ1'��}b��ȓ��}�t�� ���Ŕt��p�ȓt�(1ا�ǖ1�� �.aL���S�? �@���+(�1��.eD�L�v"O��¥�n�Hm q-D�u+�X�"O��*ޓV�I���%_,��e"O,����*Irl)"c�I���b"O�}�siy.��GAy�\)�D"O�IJ�� o��Ɂ`���Y�\M��"O��#�ׄnX�#fG×�D��"O`i�fS#)��kƃIl�u"O �I��	�j�*��A�Iz���"O�;EI?R�U0�)�+�u��"OXD��Ivo���A)�y���U"OFQ���Th)"x-iz
��� Q��y��5.��Q�_�I:��c ��yR��6 �Z�R��I�n���S����yB�%�0���(�T��2E��y��a���@�&R	i���Y�yBDQ�q� �K��5Qcv ��y��ޤW*����i-W 9�c�8�y"�H��X�"&��LHDHZ2l���yI>\�d!囔U�P��.C��ybc֎��djg"�O�n���ԛ�y�ㇵV񎰃����Kj,e�vK�y�`A2Lw��YP���#�9s&��8�y�KK�EzZ������eb�8�y�͗��]8���	��'j̆�y"��y���a4�}>1H6# ��y�拞�حc�G�% S��;1�ۜ�y2d�:`%8���֊e��⟴�y �	�ejSB�E��{Q����y�������Wn����!1�i���y���E���7�X�j�Z��\��yrs>l�(Wg�--��ĵ�y�-���(�k�n׾����4�y��ȥb<�=���6aM�lh���yR ���b�14��Z�`�g+�B�,=�8��B�=�����,9\Z�C�	�l�]Zg���_l\�1��1W��C䉪K�&%Ô�:*���A�� b��B�	 p�t�cb=�*�����GؒB�
6���:�%��J�eK0F�PC��4GC�d E�-7�����[>C�I�!�
��H�*C��(��(HiC�ɛ( �Y!tK�~ъ���ӷC��B�I1 ����SN��B��S��0�C��1{�Ct�Q�?�2�0��9��C�ɽ�R��-@�KW$����>��C�f0��&O�3p9��Q�K��~C�2C���W�����FL��B䉖�u�V#�c+��5B�}��B�I2l$��2`��eמ1zЫĨJ�B�	9x�h	�lQ�sS�=��mD50"�B�0p�|����HO�y�uk�n��C䉢hb�+'$���ʉU�ϴ.TB�:����K�>��[e@�x�B�	<8(�����
�@ˈ��V$�J�C���&p���h6: �f,�6��C��1(���[ O*\L���lG$m�B�I�Mi1zu/Z�k��)��a��BC�<�2�j$�^�4�X5a�e��B�I�hX(���M)W��JGD�:�B�	�Y���C��2G��L�6(��V$�C�I�!~4�C7~�ð$7I��B�I%�]���K�-��4� �דY��B��n���$��R�6�I��ɜ��B�)� R� �M*%���"�gY	C3֬bf"O�t�����C�T�r&S�:,�YP�"OX- E��?v|���fοbN���"O
̸֭Ο��r�K��b�~�!�"O��cF�N
?��P��� �)s"OJ�p�k
J�ĺ�a }�4�B7"ON���i�6.��:j�'J{f�b"O���Ŕ�&�H�l��@��X6;D��� dƂ;��Ţ��6�%���7D���������a0�ΐMj�x��`3D��rł�r���͌E�P%+0D����+|E��A�B��al,D�hj� [�n�-ʆ��� �>U��5D��
�F�Bʜ�#�-6aA.D���щڣ(if��C΢Pi��T�/D�X�ӕLLj��a���3"�ِo-D�tiGl	�1f(�(S�t2��7D��A�L�u$�l�W��a�b�qm(D��2T��d�4U�WjA�}.�0��*D�@�,�~X6"�d�;;\H���3D���fk]Q�	��n_�x> p�/3D�$�sn��vL%�Q�I�s�r)T�/D�H�*�C��8ڷ���p����?D�Hsѩ��Dq�� �`��Z�"D���ԢC����B��1P4��?D���`��C�4M1�jK7y��9Pg�;D�\k�.��t���!�V]�~��g�7D�@�7m݉���6B� F0J�b6D� ˶&JEa�pQ&��_�.����4D����
0�|���ឞ}{���o?D���&�N'ʈ���l�@���>D�SS����#ٕb�B�H�>D���q�0(W�P�-Z�U��/(D��
&jџ+�u�)�.;���6`'D�K�������#��(�bL D����+K^T��M�&*��A�g"D� ��?=�*\1'D�z%���m5D�4��>->^�p�E�4Sq�c*4D����2Vlf�)2����W�2D��BE��NW���@쁓I���C�-D�\��&γ$�V�ږ�y#���+D��`��<s�������n��m3�Of�Y�$qJ�˄���$d�b�������M	F}��/A]Z=Psc/D��*�W5	B�hg��Z �b9D������Fڔ���A�,?M�]��6D�����_4c���kF�)�vŹA�2D��x���"b� Kp���,�he#�!2D��a���K��y���í�xY;P�/D���vC��&g��s�!�5G~V�k�;D���T��6���� �s�*U���<D���@��� �`a�!��J�q�S�:D��3JG�d'<�ME}� �
�h8D�����Y��=��HQ�`2���6�7D�T��[�
zɒ�7s��Y�$5D�h[�aǿD�@J�O²(�<���6D�{R���p{nT	�& ����@6D��q���ʆ���]�� mr�"1D�D�c^�$ajٹ�Z /~:[!:D��ZBl�	���A��2�V�P�5D�b�j�5���� �ɐZ0&l16�3D�ܚ�)vD�Q1��<Od���G,D�l�C˖0i��X�{�Rt�S�7D����)Rܼ4bR��K^�+G�8D��  A�$�#�l�Z�f ,��x
"O ��ِIRp�hM�M1�(��'3�����=M�Դ��c@��9�'���K����]��<p) E�'t��Х~��R#��>8��a�'��Mڷ&�N��ؑ��uBx��'�<{�%A�iu�Q��P�l����'��s�%��8��]����k^T�
�'�.U� �p̙�Dd�=c:i
�'����S�\f�$@b���'7�m�u��:Ut�)��G�g�Е�'^������=R��X*�$���'W*�[�ǃ%C+�����5��K�'M�`Ѓ9'2��y�n�&�R�'�����PZ�E&F"j`�!!
�'22�"�m��P���$_�|�	�'Z�$�P�P�p�$�KD�D3Gк-��'����Ҏ �-�|d"93J�)�'@N���@O%F8H#��+%@de�'�Y��Y�<�й��kL U��B.Y��C�#K{����bG�T�ȓ6;ڜ'�`�ȤO�#@��І�U��jg,�A�d�%a�w�8��ȓ&���5�ѻ�|�t�ϹAژ��ȓ�:)�f㖁'F< q2��ko����S)�U��d��u5fxJC�X X�4C�	3T)���"'˂R�`���	�2��B�	�	�m(�ȑZ0|Y�G�i�4B�	�X�RE���AP(�|W2B�	u*�
�U5�l����=B�Ɍ"ɰ�A�*_�q0���T��C�	�N���1���7��1���)��B�=C1�i���.�H��rdԶ�B䉖p�=`��gG�T{#�֔xJ�C䉈v0�$`�$Yc�D�a,��2�B䉿JӠ�І
KrL�4A��v�zB�I�`/�b�E�*:fV��?��{�"O��P�ަ����GBP01�F���"OR����(X6L����vo��X7"O�=�WM����S���qg-�"O~��BP;'.�M�F�%yOJ�g"OB��t����=���*=(�f"O��T�I��h��5
�ġ��"O4Q�V�]�z~����ڭn��z5"O��̶��(g͜�W���� "O�!���%l
�5(�Aȏh� !!g"O~XzB��' ���C�'��� "OY�,�J��ЂV�ŜR�<e��"Oԩ
���}/&�qB`�/Zy�W"OFdj3	�g%  .L/S$�dɀ"OP�2�D�yiHzӯʫ'��c�"Ot�'(
)h��2ϐ9
� ��"O��:��³u�z6�ڐz���"O��!�A�4�T�
��y���3"O�0a��� 9��I:��Ǫ[� q"O��׌��V7�3AjǸ�����"On�f�[8?�⁫�D3PY>�`"O��I#�AiR��*�&~hf��"Ov�)�-��Xd#dS6SM
]("OT5	0�X�v(�D��.K7^��"O,9B�"��L�H�m�\3|	��"O�p���W�kax ��ο?3���e"O��K�e��1B�����;+�ta"O���2�	9F�
�;�h��\��0y""O� B�R�
܁l�P�ٶƇ�H�ށhg"Oh��W$9�}
�Bo�BT�"O�P�@(4�>\����%{4�5X�"O��`CD_:e���tGԞR,�ju"O�@�'�=թPGI�$qk�"O����-]�R�8�F a�I �"O6y1f�I
A+2���N�J@'"O�!�%Cm00cE>G�4��"O�%ZB�¬mqz,: �Sm2�'"OL��e�Z
C� 9���J��v�s�"Ol�����^��0�hZ�}�.�z�"O�U
����4PҨ�	]��� t"O��4G�U�\ s.���tsE"Or��d��2��MU�n�����"O����DҶ,'�Y�'��QE����"O��#"�PnZ���Bڇ,�,X�"O2 �2�ܚ�:H�����4~!Z�"Oh�ʔD�
�Fp�T�8��"O�vϝ� @��U�0u,��t"ORV�U�` g&�����"O�ŐCI��4ґ�
8q����"O��@MɁ���(�bɴb�j���"OV��֠�zWl��C��!,:�$�""O�$��m�kH��g��	+(���"OҨk1i��j��d$�Q&tY8T"OL�qv�D�W�:���!2 �"O&��ŤF*Y�l�2������"O��Q�q-��3�mB��d�"OZ�r�� �
Dn�5x>^1�"O��2�L�F���r��10H�)W"O��4���T�N��E�߈/9<�R�"O�)i4aA�+���@���-��;�"O� �F.�:E6�̘�b��  ��a"O�`�����P�8u`OA�T*�)�"O�iD�Q�w8�ʡ�C�L�b��"Of�W�^:6"z�3@�6P���k�"O���� �2�X`��.���"O��!r�N�l)h$�?m#�qY4"O^���ɀ:n�`��''�,#�p��"O`	�"��9ڄYA�аVV���R"O�,QC޶X�`YSu�ã]Z�ū�"O�ݒ㢀�<>:�����yK���"O��ч^����s�ػPFl��u"O`q�$�L"����/40HR�"O������>ى���&,��"O���dіd��u��K���2"O�"�B� TP���s��y��X�"O }���']>�bE��g���[�"O&|����p��}�s#H�dy��9"O�Q��I�azh�W�I�yxn�H�"O�-HҠ.2�IЗ�P�1U�eї"O�ٸUg�38D<daPA\���"O ���3L�(��X!|���;u"O��ӗa(�����3pT���1"O��rE���z����A�ieԌy&"O�����ϫz�8�#�O[ Z��R"O
�;W�$�5+5/O�"I��"O8k���4(7�ذiZR�0�"O��"�͓!SSB��E+�<%:��"O> ��A�B�ld*E���͚c"O.Ɋ�����I�G�@5(:��"O�#��*�
 �P&؞t#^���"O\x�t���{��V	5~*���"OR��ß)6�8�qs�ZMd�Ч"O� ̥R)T�Ĩ��H� Z�BQ"O�H�&��`$�b2���Rf�02"O�=�B�`�����`D�,Lx��"O��k� ��ȱ�O�h����u"O��pa`O0/�>�+EoV�iۀ �"Of�d�j�en�x��,�"O�SS�΃[j�Z$@�!4�V�b�"O���B�)Xp�wN3 � e"O����h�=�ڵ`3-�;� �ir"OLԸ �"�|=g���=��U"�"O�y�c	���r�OX-<yj��t"O�Z"$EI�X1q�C�,V���"OkV~M��L�1Umj��u"O��q7E��s[j@�0D�/^b��"Oz�r5L�aZ�ax��^2�6Q�t"O:ĠLO�����#�(�K�"O�P֍��[��|�@�P1���J�"Oڱ�1K��b�
�N@�VT��C5"O�rDX�rX�����^6XB�"O��K�m�_�
�P�mM)7�츂"O�I��.���$ ЌW�~, �� "On�Id��u�\��K�:F,L��""ON�c��O�9ZH��)Y:C~"ܪ�"Oз�J�OĪ��y,"O��6��.t|�yQiE�?�t="O�5�4-�~��əg�Qm~X��"O�!{�h�C��Um��LTn�q3"O�u�r�� �VX5Nۦn7�8"O���ޢإSE$d ����"O6@yƩA�?�����P�%�:�r�"O��#�m�X��,1%A^�Na�"O�л���N�n	�c�0a`���"Oj�"��&}Nʨ9����c�64g"O��ug�\�9��Ƞ<�L�"O�a� ϟC�.���٩K�д��"O��PǗ)V���膱9id0"�"O�8Ȥd�(�`"��
�B{��b#"O���a�	!Y��s&FGPn�ق"O5Ʌ�Q<?m�9r�OH��0�"Op�Yt�=`�,�D�s��X�Q"Op�1/�<��c���2�a�"O�h{��
V�HT�`�41�1�"OE�]/6�G���S�"OV; n��k7h9�u/��4СX�"OFI�%O��HӺ 0�B�a�X�"O�W�A�ƭg�֐��"O�$�G�ī7�L��0�
���X�"O�f	�OL��ʒHF�JPN�
�"OP���Q�+�Z���gO�.*�83�"O ���_6,��ǲt��e"OĠ� �O*K�fX1^d4�S"O @�7mЯ�Dl�eĞ>����7"O a�Uf �dq>�O3�� �@"OQB+��s�b�{a�P���W!��= ��YibL�O�����K��VQ!�D�K���rf*R%Q<�KU��<l�!�Tj�MJ� ����JT�ŧ�!��^F�`�b놃d>6=i,K(�!�ą�dZ���^\<�y���V�:�!�W0U0R���,7Q#���⇣N�!�I!5�T�e(!<��� }:!�j5:�"'_ r����ǁX�9!�$
=f�,h�b�?k�DhJ㢞i!�dǹ��dxUD������ʻQ!�� 2]�q�I�969��l��P#28r�"O���G�h�@�5��Ό�uB%D���t�S�f���q�]����j$D�,�NG04����jW/Bɐ(�A�"D�4�t��9�fp3����^EP ��+"D�hHc�U5_d�;"��?]:�0�?D��9�ӵyJ�c��@%"�°&?D���Ե%�<}$k��,�0�a��*D���Ab�X枱��!ш0���'D��ʖȅ������O0u¬�Y�;D�����(P z4#�"4|�~���A9D�� ���=?�!� E
>+NzI�C�5D��Q�k��d����(
4(	�k�g4D���J��&�0�r�b ��as(D�hؠG�F@�0��A� ��Ae%D�,b��B�D!0 
 k2�@e�0D�$a ��0Ƃ ����!��$��g;D�(��6[�z��W'F�z>B�H&":D�x�IԬ���Ҧ�1v�C��9D�̘��m��D�Nޮ@��8D�ૅd�:�b�䯀�n5���׌6D���,W�|�X�k��B�V���2ů4D���voU�-i��AD��&~�\�A�&D�D�T��9m�}��G
F�� D� 0(Fm�� ƨW�d�(� 1D�(����E��@1c�I�x�8�)9D��K2m2n"]�"�u�@	8�8D��Fォdt�$�+���K%�8D����!��v���/��x�t
5D��Q�.B�%�(�r҆ %'�!�D��dAF�P�l�����rgf�Jm!�$N�T����l�$2Z�;�J�=GF!�$�F'x@�4A��a�b�"�I��$!��	2��=@v�� 48�hI:�!��ט2��"�#�Ni敺CȌ��!��ߥ��ՠ�+N�|YF���P�!�$�*S�0P32��pa$,�#n��u�!�ěa��B��y��P�U!k4!�ċ%�>����90�1���-!��Hx$5�`�c>!�$W�f�|0��׮���e��	(!�d�4q(�A�uB��(�P���"j!���?l�I:�Z�,�0��H�!�DH<p9�\j�����&@ϳ`!�DJ8��Y-1c��ӍI�u|a�'b���a�2LX��d�j�
1 �'̀�����S���83I��_Ǻ�`
�'ն�q�����)��g�^Q�q��'}���C�C�`�$hDA�C����'���рN��7t����=Z���'�*�S(�$Na�Æè�j���'\���#M>r�񃳢�39 P;�'�v�{_P���s$@W#`�x��'H��i��3��X�#���&$��'�:�rp/G�dLX�sc����a1�'Uࠁw�h��"���l��'���{ƣÂ�\�2l�=��E��'�㥭O\b�B.�R=��'/�C����h� "B' �0�'���oD;`��9��
�'I~隕Aҙ[X���A�נE>niS
�'
����8���[a�����	�'����F�7�JD�3mė}/h�(�'�Fi�q�D�� �E,	)������ ځ�/ґAt�s�c�Wz�۔"O�b�E@'@�pr5b��ʖ���"O>�wI��\����@��OS"]��"O~��#b��6]�0�H��,�x�� "O9X@f�1��p��&[0D�0����4S���$j���'���X?�r$ŋ�?ӂ��J�Q�6M!`��.=O�8q���?��
Ą`�0"�7��, .�V�6��.k>�P���3A�h�SH��
�X�m%�OB���a�ԺA؄Q`"�s�<�UDH�7\����|?�Aqf��d������'!R� ���?��d�ic.�TLD9���W��h�0F�O��O����O�p��늑8E*��5`�8V�P(A��'�7��O<6����b�� o�'�t���Iı'N�9�I9V]��0ڴ�?����?��'gS��p��?q�4��PID�!e����j��a 蘩5����(1�$��Q	<�֥�'�����X>μI�t�ӌ >
Q�'	�)e�7��/Q�P雐f9�"$QgcA�FoB��;�u�F)���ḧc���>&q)�!P8H,�@�iuH�����?9�O�T�sӆe�O� �؝��E�(4p��O��%�O~� ��8H�$U��h�K��<SW헱osfb����4�?��t�i�~�S��/b���G��:j@1�O����>
�+�C�O>���O0�$�������M3�(+��i�j@	{ ���lG�g��A����� a��ނK���0��O�� Dx���6p¼YD��8դ���h�y�ڸ.ua���MÅz�r�s�b�a��B}��6�TS�$��~a��C���f�c�؃7,��3V|���ȟDyI<�-���g��;�T�I6R��A[,��0�)�矠��NL6� Z��R�p�1�P���r�ҒO�ퟶʓc����2N�jI`l��� ��8@U���*a*� ��?���?	�G͍�?q���?I��:�M���YN�8V�.fp!�f��#������X ��I���Y�'A�}��f��~�P	n��Ȃf�6I�9S�*Vw�yu-��<z7�e��}�?i��Y���l�G�J%h�ꐤU$y��dx0!zǽil2Z��ã	�s�ӺӜO�v]�� �8����Ċr|�5Q	�'�>%B'N���e;`*�6c<L���'�66m����'�J���hb�H�D�O2�'#@x�K���V�(3F���X�0B+T5	��'�b ��ؚ�H�Ɛn|��Oқbnj��'+�t��ٝ3o\��_�a�d Dz'�	Vl���V

vp��۰@]�֝�N\d՛ i^�W��[�L0�$���[`��&������N|��4�5 �E_�3���j��ML���'L�O?��� g��� �ѕ.�ZI�#aE�@иD{���nj��'$��ݢ�+�*w�E ���J����?��3GX� ��r�t!��3(�'���n��`Y�,�������`����V�4��C�+�tZqK�,Ay�@h�I^����P>=���CIX�+b��lĵ���3�����@�A�H��Ɵ"Or�%	�%_��u׾�N]%?�ضe�D�3ͅ�s�=T��<�<7m׈yu��'>�6�O�#~nڈ+���E�&(
�er��c���I� �?��d{"ꁻ�)�?��(��jK%�Q����4�6��`���H�?b�"�r�ʣ~�M��#׾���=	�eT   �   ]   Ĵ���	��Z�Zv)Ċ;R��(3��H�ݴ���qe�H~-�8L,<���i�n�?
.Q�0�đmz(�Ӥ�._6��)�4<�>��' ��0O��@6�ʖ���:"m�&To�pS�Y2j��RߴZBqOR����D^*�MW�[	A�Ʃ+oY�Y��,���V���D 8Qf}I�4$���.�응e�:ל�;R}��c��e�Hu�Ҏ��K$ ����6)<��'���v�Z&(%�OR�2d��v�4�
��ȜJ���ʡ��g��o�$�?i�'Ed���=Q�)-O,��U'J�D��\c�(y�S菳tT,hĭG�WĂ)�O>��M8�zrF�O�mےl�&�,a�fg� M-BA<O��������OH�h2CS"g(�\�-�A��$�r�p�'��IExbkN}�)�?-|���!�T'.��Q�L���W��3F�D� )�����%ߖSjՙ��ʈ.
��J�A�'|ZuDxR���3�|PS�C�����tf6yӨm�}rBK�'�N4䧭<�rME�{�X`�b�,v~�l(O��9��D�<��'}l8�Q�20*i���5g� \A"�V~�'�%Ex��Vߟ�	wA̙D���1!.��8n��X!.&�I�8��x��x����w4����4zxӤ�\.�~R��x�'��(Eyr.ԱtCDI�s�M'�`R���?i$�d}B�8����t��u7:���*eB��t� GOR(�P�H�ƇN�7D,�O�%���\�'}����C]~��t#��� g͌�	4��M>�d�ۈ*6�Q�<�I�)�Xa�(Y�=lT�fЯ�PX��'Nl��@ ��"O��Y�N-W*`���R	Hܩ�D"O��h�f�;P�&�@2�"x�a�3O��x��� K�JQ���ʤl������f���D�4�O�jR'�j�V(�l�P�.��u�	�]�9r��B�T��O:���b�F�44X�(v U����'Q�����3!pĸ��EY�N��I��O��C&��,��l�m
T>��¦��@t�r�lF>]���pH5D��"�/[(j��	���Ĳ���YRL�/O،hVc��9:`<%>c��;��&���į�%!Fb1�-'�O���פ��]i�]k�f�:�%KPN"�í2���B�'�~}i!`�'j[+��I&A�����)��X�KY[���O�q)T�ڱD�� s-�E��-��'aL��⊯\�-3%�>�fix�Ox�Ұ�X�/��If�[>a�    �    R  �  �  &&  x'   Ĵ���	����Z�/C�'ll\�0�|r�'a�	�Dط8��0b�
�<�}#�'�t4��B�h�dt,�:?������i"x�	�-��K����1Bʚ�HH�� Ҕz�J�[�.�0�|)`��u䨉:�Œ�_2Ii�$]�-��s�	��	-�i�V���LX��92��6�x)����sA�)(E&X�9צ��
����q�`˯do���ЂL99}�4y2�E�C����>��(J�"���U�i�����m�<�e���Vk�$�r���3�,���E^�<�Ѝ3?�0���x"���,�]�<�BcQ�P�nЈ�"R�	cT����M�<YDc�r��1��Y�����F�<Q�ձP�҅����*
8�P{6�B�<鲆
(z8���J�%~A�C�N_�<1�!+��|�p!O!gƖkB�F�<��o	�;��B��[;Q�xYq��~�<�և�+}xe薋���b��d�Qf�<�!��.0� �a�=5l���
d�<��"Ι%yMX$(��^W$���|�<I$l[?E~*�l�!Ha�T�C�y4xF~8i�bL�qȂp���y�)�	{O�|���
�txf���J�ym �}Y�*#*��7\�@V$C7�y�M+,:Ѐ�JB�9�0C�gN�y(�q�:�$�M⧄VG!�T'!w���3�X,B���]!�LJ�.h�wD	�6�a�P��(v(!�D4 ���H�o"ʁY��ѻt�!�$!W[V��1΀! 1��F_Z�!��T�Ms�@�/��j���wFòk�!��D��(��&o��B�/E�!��q�%��O�2�&yz�΅�k�!�D��6��<	o�R�(�`�M�<!�ĜRq���Wc&V��K�-<!��yy�����b$�Њ�t/!��H�fؠ���0�����V9!�C�p}܈r�j��Se<���Α�B䉭W����KD��	 �3|pC�"Oh�q[�	 �j�h]j5�փO-�C�I�"�� �S������0��C䉴([4��BH
C��]�2���1˨C�I�3��c0�N�j��q��&����C�ɸ���[2��1-�Q&�̧:�bB�I.t*�]�7+W(8C�[�/Р"�2B�I�r�@�D ���H2���
B�UCL�⋀2:*�b�;|�C�IRU@��m�	8���k��M�BB�	/���ck�u���"D��!:�C�	8W%����o c~�E�D�î�C��
=�x�0�E��-"0�ˆ��7D�fB�	�+���ħ�bm�V�D�y�hB�I;=���+� >�@�1/�4+%XB�	�~0��ԧ�3[i.i�0(��sxB�I,\ ���d�ѵ3!b���S�BB��9�0H��� C'��Bh��)�C�I\���ao� �Ď���C�	;A�d5`���/}����C�(%�C�ɯmh|dZpe��o��0��-�eA�C�	��f����N�h�\�'F�B��C�ɣ;���{LG�s�r�
fσ�l(hB�I�v!��đ$8)F��� �Ju8B�ɣ�dX�g$�6%"��P�S�&Z�C�	��PE�e3}�]�g"ݯ~��C�I>�a��"�1zr6���"X3ZB�I!^0���"#�-<����DX�L�B䉛jwL��JݳM]�X%��`8nC�)� RL�6g\�F�
��f�%Z�"OmQ�2����w	I.80��"O����,���"��c�N�3"O�U��M�B��L�sȞ�M_r���"O��V�>n�A�l&X]+q"Ox In�>�j���	��v�lA@"O��Ct��C�����4E�f�+E"O��1�ED/Cb4�����`)1�"O(� ��bR�@��0���1"O��1BոL�|<"<H�Hq� "O�k��&S<EQ��-���%"O� AqВZ�RP�%����S�"O���cLa6���\Ȉc"OJ0� &Q�z��@I��[�_|��"O��V���:C�t��GB�U�p�i�"Oͨ�k�7���s'��1�U[a"Ov�+v-N3�j@��e�[ߚl� "OZ�b/2�tC1�M�dȞE�r"O8��O�#3�)YE�R5`|�e"Op�ʖA���8�f	�}���"OB�xT�L�P�a��7�%!�"O�8ش��)��t��닦,c�}�3"O�)��M͜�� ��JկZ]�3"O(���	�*�\XtI�xJx��s"O�Y[&�K�AT%���E����"O�-��-Q0 ���K@Kۨ\{XS�"ON9�F�'Tࢯʿ;Q$��"O|Uc؋e$�r� � V��}��"OHp�)��.�a�
�%O�� "OH���DG
�B4�q�L?D�<�*�"OJ���
.q�u
�9�>�s"O�K�%\,NHw	ή8����"O6�˗�SfT����/
��h��"OR5�A,!L2��OS1s��3D"O>q�&I�D2��bNح)���%"O��F��1&ʄ�#��t�#q"OX�����IZP�����3�X��"O^�U��ZrΔ��D���"OL�auGH�|�P+�Ů���"O
���Z3R����鑘b%Ъ�"O���*��? �	�hcܬ��"O�{U�;ø$�ceH�e.���"O�)��ٵj�����Q3'V�@�6"O��Ң$B�O��X�j�ܑ�S"O�Ds���4��R�hN�C��D�G"O��U�O
.1���SD�2��"O�$�R�?OH$q6/ҹ~0H0��"O"�SGF\=RY�#�A&�;�"O,hRe��9Lv�]�%�������"O\�s�M�W��	1��)�BP:'"O
y��D��-$�S�0e��Xxc"O��"�'I�pZ~=2�N�:�6(�e"O�1�7Y�i�PO��85����"O�)��͂&�ikw͕9#�2	�r"O���@�R�������'�,�i�"O8ɱa�٣g��U(sA@�t��e��"O2��SƐ(/9�]ЕG��I� 4�"O ��5������&K�h��\�v"OdiD��"y:�3�>*�"O\�K1�H�]
���
:<�P �"O��X��3�f!CvkFq�d[�"OD������RA^��ֈ$�"O������B���sf�G䨚�"O���Q�Y�8�
�{`�϶X1��ڀ"O� <�G�S/N��0��3M�,�R"O�T%*��x�V!z���|��"O�$r�)��=�l�j���
0�2L�A"O8���I�hV��  ���0�.�c"OT9rn��.�{h��e����"Oe�&o�$t*8Y1�9b��"�"Ot���6���b���bVb�XG*Of���̌����h�H��m����'9:ٚ���-�T� ���P���'�hiC�����K�^0�	 �'�>�bH��^�։8`���R�v=��'��5C���t� �:�ڶi�'��@feC,Sf�P���6F� ԋ�'�t�jb凌0��=Yu��Ky��
�'�pB����<4�$	�,O�Y �'P��c�a�7u�,��ۋ
!F��'Z.@3拌5gf%xg/ܟ h1��'�}y�)Z�=$!r�E�A�4�p�'��xx��o�& ���(w���0	�'ђ]yA`�)"N��"���Z�Ν
�'Q�������!��O�_�* ��'����a&N�{���ѷBR�<�'�@�0�c��,#PQ�4,̋L�x=�'�(J ̊�.�@[�`��~X�`	�'�d=`2��R	�mkƃ��w�+�'��� 針ϊ��1�OOTC�'�6�pED[�.�bp�ƌ�X2]�
�'� Yi�%;
*��E�/_k���'�hu�Ǭ	!f��,��a�G��\�
�'Z�T��x���U��͉�'H��#����xИ$�U_	L� �'�z J�*�&j7�ˤ@�6W��;	�' 
u�E��& ����"Ҍ]	z-��'TDQ{�!��_ H��9b�8�'�Xbc	4qw����!�Ϩ��'� �CmK�o�`��g����A��'��)(Eg?z��-�!˻5��mQ�'�<��Gˋ�[�H`��З7'�t�	�'��Hr��33Z�J�a�>#���P
�'@|	H�i2yN�@b@��1�	
�'�B��e�{�vlx������'�a�v!�+�Is�̝�Y
�'��djG� }��Y��K��3�'�v)�!i� 0��́r��$t��	�'L2���B��(�`'� � �"�'ir@�*M<nh��+Q��F` �'�nL�A')���ĉH?����'�d�`�"˘?+�� �h��<���
�'��q0��Ǣ\f���7���3Ϭ`�
�'�f�[���(U��`����#�$[
�'(̪�E�.\ԡ�1
L���j�'~E�s(*�ԋ���O�f���'��yp N�%f�ơ8$�ͧo�`"�'�49�i_���E䋘�8)����']�u{�l� �*�ɠ�3>1��'c4 v��@�T�JC�:�X�B�'� ��K�/��)�s�*9�\�	�'�$�
E`��1�tAYC��(t�	�'�0�j�D#H�<�ӌ/)��tY	�'4�C,O�=�<�g+׊5/���'4)ˁ��,։H��5�`���'X�4���X
G���iB*�o����'>��r�֊.���u����5!�'�A�(ON����NJˤ�+��� ��H��"4	�	۸rb��t"O9iE^�U<Mp֯ϲ=��� `"O�\�v ��0��E�3��\�"80�"OVI�
[�8p6MYG*�<X���"O�a#�+�o�H���F��Q"O+M��l4́1fO��{��W��!���:B���H�"A�ls��ޮ�!��T��*1�	D(y�(e�!���7 ������ß"c(���ʝ�;�L|�Z�����	�U���A0f��M���z�AS5}߈C�ɨ_��y��$��諤�;GO�B�I`�l�s@�"i��C��B�Ɉc]NL	�Y<,p>��B͍!_ B�I�"(����;�J�*ׯʈt��C�I�'q0҇KL�k�Dl�%���7%�C�ɘa6x(f-T��!I�R�JTB�	�no����N<J_ar�D��$)�C�I�~��D��A�$9X�H�3:�(C䉛62l�����:Qs���2A]t8C��
�QČ�uH�m�����4C�ɰ4,�9��/�}�DS��8HC�I:s*�$sB��}��M��	۬<XB��	) l�
�ϗ <TԽʁ�ܝ�\C�ɰw�,02��"M�dq-�#qC�I%A�4��2��=���a��U�[l2C�	kS�"ң?D�9�%�&V�C��#W�
e�aS=)R`�	`�`,(C��
����c�@9H7�1��+�L��B�	�7�V4��KD%���₢͇*��B��pT\���7bJIR5Ν,U��B�ɃG��8�3�WvP�ȳǫ�u�ZC��C�va�pIW6IfX�Y��G���B�ɯ�
���N�:J2&Ѐo�r\�B�I�Y�d����<#d��$�8D�\C䉾7ܴLRG�§:MrӧN�q)^C�I�>e �b,ؘld���a9U�B�I1>�,��<��T�eFL��~B�	��ؘd��l����i˅�xB�ɯwc``BƊ�9j�p�� ��>��C�2do�X�B���d4�u�˙nK*B��#Q��E�E�V�A)<*��\�g�(B䉁R��� iؿ6�+fě4B�B�$\�� ���҃B����M3�C�	L�f�2v!˙{+*����6{&�C��'^������U>Č:a�ȵ{
�C�ɹy`Jpɒ��	d׆��0��2x�C�2w@v�CƬ�-�\�+�f��D��C�0b��a��ϑ4���`�	y/�C��h��b�A9`���;ׂ_&"�LB�ɖ`���p��^33<xu㥍><�&B�	��Eb�J.z�H��h	�y��C�)2�H��L�Go�Q��JC
M�C��<C����E��N ���l��C�	�\<N��#�G�9�n�!���[��C��2w@L\9p'�!&n:�t@�t�C�ɸ�0���H� �5�h ��"O�1i��$a1�%��N#���w"O��။�=�;�N�dnI��"O4��1cM�{jY;��@�~4�[�"O����+U2�>Ds�,1�(�D"O�,��d,
� �LU�e�h��"Or�X7��'�Th�����Ф�e"O��
��ݫ*|�!�*_�{p��"OV���mځ-(Ah���fĭ9�"O� ��Au��!pe�r�#VmC�m�"O��B&D��qQd#)�졐P"O>�&���T�
	�b^t��E	�"O�������l��YG�&���"Ovѓ1IZ�~�B���<���"Or\�Ԉ��Q8��Ǌ!;�"�Ѓ"OL��"A��^�|���}�̴��"O�(��*ٵ5Ȳ]���="1�5"O���#Ip�Q2��E�1�"O�Yk�d��CtCƣ�tzd"O�B���:�d��vǏ��~�"O^�h��!�0�r�EQA�|ZT"O�e�b�Z�E�X�7ś�0�v�;�"O���קÇ ���c4��3	nd�H2"OA���D:]�:�+�dC�WevВ�"O��鐀љS�&�1vAD�j>pd�w"O�Ѱ7O����V�X#���%"O�|�$j�{[`��$��K�80�'"O��c4&ǆuw��'B� j����"ON=�/B�H�ോb� M�1[g"Or�
e���ޕzf���5�
ŨT"O���g ���}�a��6���[�"OB�Z>]����ɋo&lA5"O��2�.ɥ"��E�'��8&�H"O
�O�!|1�$���5W�8S�"O���皅t��p!	K�����"O�(���L}����+D��}h�"Oj`"��
�4YR�VO�"J��"OF]�f'J�~{���Q��-j��"O �#$jJ�& �1t,D�o_��(�"O�$��Z� �:�+��$<:�S"O��Z��7"M �2�X����"O�0rfhR;j��T FfE,�� pt"O<Ձq�٣<a��Җe��|��)8�"O�Q`i��~�˳N�M��E��"O�X��]!j�z�ʲg�$���"O�RQ���:x@�&旯Mΐ�%"Oh83���u���@��1r�b�+�"OBU�&e	�Wr�c5��rߊ%�d"O�[V%�	�00���NΞQ�"O�Ѳ3o[a�D��?mZ�*f"O$�V��/?j�A5BO�gNr�a�"O�Uk�e�xz��O�6C�I#�"O�����״��狊�ba)�q"O�����r8�r��5X����"O����Ώ�*dX�RIƀ@T��`1"O@R�+cq~Sw�֨_>�i�"O�ɘ D	T@��� ̯Tŀ�		�'�J8�Fo_;iQ��HS
�b9�'A*���+�
Z*�S� ��>�+�'�:�u�
~j���rg��	ޤ�'�"�b��$KU,t@��M3���'��8�H��dK��Q1�^~
@��'�hh��Ȃ���yc�ȶ�nL��'�(���8�ԅkU��x���K�'�P8��
LAk���.��h��`!�'��j��^+q����dgN^�4�8�'`�A���{��e񠝉P��h�'=b����b��%
Q�]�LRFD��'���Z&�@G(TK���G� �
�'�|�����<�8� #�P�r���'���5� [�p�oQ
	?Ҩ��'��iD�������E��t��'���hAe�0{A�]�@!��s�"O� ��it�̮w�X#��U�i���p'"O<���F]�h�H����E�)�
#�"O�H2�� &�~ŃW%I�i��8��"Oּ�Q~AZ��A]��M{�"O2`����;�e���<?v&��"Oq@
,0�H���9���r#"Op���h�R��%͜A�X�4"O�bdm��.�n :��¥w|N	sa"Oȅ����~8ȡA1��q�A��"O��S�R�@Ъ�����! X��I�"O�u� �0f�Z=�ꗆe�
pb"O���G&ɶc;���J��t��<��"O�Q�ggd\��(ң=�zm�"OL1���>V���Є�D�bΦpa"O�lS�m��?����W�`�
��"OPy��7	r,P���"�xʆ"O`�������X�=��Y��"OT�ڥ"�*\xi�� g{�,+c"OP�Pq�C�F.6�Z'��^���i'"O�����<O��Ex&�Z�Cy(U˅"O������z��鳒�!<O`�Q"ON���O'Fp����Ȥ[6�-XP"OJ0ˁb�>(��ظE)��T��U��"O�Ȁ�+��*�*%ZI��w���R"O�	
���R��D������c�"O���!ڸ��q*�ǋ�`����"O�䂐�@z�܌���K#����"O0��"��(Ј�j0-º� T"Obh�r�.+�0C����,E�̹q"O�S���|ء�&�$=�}X "O��R�?��[a`��/:� �"O<�;� �=��4�q�_�&��"O�XǤT�t�\A9E�ǒy�혰"O���N� /�0IA%G�u�Yv"O*c�&�t���r�B�T	� �"Oe��!�$9t��f�_�"�|���"OR`rv#LHH�I�i�4B�pLQu"Oڽ���� ^��E	�~�p��"O��AG
�>�>d��g��� �"OB����[�P��d� fU �=�"ONI,,��"Q�**a�*[�!�d�7:�d�V�Q�~�6����T�D�!�Z�A�ܵ��m�	E�bO��!�d��l2��#+�2 :�`��� �!���46(���J&P�y����	W�!��P�o�vMZ�B�|��1���!�C>^�X���{��=��얖o�!�ă�<ۼ�2f���I0=�JD�e!���(A�^� 2�Z�F�l�K��A��!��;wA�\�ש,H�� b�@5!�ϓ(����m�09�P`˽q!�D@�Gl���]�O��`g�1m�!���r5a%+°L{��1�Ơz�!�D
�;@X���N,�[���Q!�$O��$����b�ڠGX�,a!�f� ��X�~_�mA&@�$!�D���l5�#�JW���q���>!��/zV��I��mSԂլ��u!��^�rh����=q��sDMZ�Z�!��5Rz"@�����6DJ�Z
&�!�Ԅ8j  �d'�4D���F�!�$];��!4M�p���Sc�V$G�!����5A&O�R)>=q0$�!�d�6tF�cB�;r�Yc��j!�� �$c D�u�ʌ@�R�5/f�s"ObP�����C"��:P���*�0�`�"O�9�J��:�H�;��&U�
5�P"O���^XI�����9��"O��X&�֕F]�Dm��`=�"O�ŲEK�6=a~ɲ���!J�{�"O4\ɒ��-+V!��%g�#"O�%c�Òr di�Hج<|��"O�� �鄌uܘ�'��O�|�"O�t�/�R<p8���9�@��"O��QV�D�*>�h���"����"O�|Cq
�1�t��$i	(P�zM�2"O��Ы��)�q�Gǉ�SbF��"OB���  �   j   Ĵ���	��Z�RV)Ǒ7>��(3��H��R�
O�ظ2a$?����H�49a��i��I��i� ]�=����V`�6̀��9X�4Z���a�'[�V��p�4�I�8QP�Z�d��V}@����2Sd#<G�5x�67�]�|mN![g
��{� < gÌ,%���`8����2��L�OUrQ��_�qJ��'h�As&N���3�f�p4�+��5��L�?{�L%�z#
1;w�Z�.���ԟ6��6D�	2K�*ְ���qn<!(��C�+R!" �O�� �%�W`6�h�X�����<���� D�>b x�֍_�Ԓ�-[�2$R��'׮���d	@�'���'�)��N�6"� mԈv,�4rhe��i��I"5��H�/X)c7�!B-�2N$K' 8�O���Ď#��� [��e�@X1$s�����L)tg�H#<��6�Iƒ�l�D�<\:��iМ�B��i�qDx�k�L�'�t�dW5@eĸ3ڳ<=��IY��'pz�Ex�p~�JÝi!��p�A�Q4��[5�ի��$�'�O������,-d�FB��L�2�H��خ7�4Ex���f�'D�!�I#e����0fZ ���C�6h$�b�( G�I�'{0�PrNЀv�(0pC�D�441�'}HDx���I8[���fKG?�d��fc��e���T�ۚ,>� �%o��Y+ߴRk�|CCJG�'t��*����u��ߢ&XTx�@�ڈI�DX۔
�^qORl���[
����X��ǈa� �:Ή�7�P��%X6�q'����(O<U��ҳf����Ϩ(2���"O,���  ��]�\	.#�p�A*��Ɇ4`�(�b�V����hR��LmJ��B�&��G=�¡:Wid�E�CF"t�p�җ#�3u�	���M��$@# �<��h
93Q�����-A"Kc�\�"�O��0«?D�0�k�%k�r��"T�]v�ʀL�<��'�B�0gTd
̀1႕19J"ܮj�FDB�'m���@��|ɠmҋV&X��דj�2i��)b��;����F�H��3?e{�N��2W��# b�Gٹ_�<A��cy���3�j��M(����$���	�� �=��$ ̐P��gR!:��I""�L|�#h�29�B䕴f�y��_�C:9��#���?Q�HA*1��J�\?��,p�e�����4����ݲ�(O�t��S��,
�8    �    R  �  �  &&  x'   Ĵ���	����Z�/C�'ll\�0�|r�'a�	�Dط8��0b�
�<�}#�'�t4��B�h�dt,�:?������i"x�	�-��K����1Bʚ�HH�� Ҕz�J�[�.�0�|)`��u䨉:�Œ�_2Ii�$]�-��s�	��	-�i�V���LX��92��6�x)����sA�)(E&X�9צ��
����q�`˯do���ЂL99}�4y2�E�C����>��(J�"���U�i�����m�<�e���Vk�$�r���3�,���E^�<�Ѝ3?�0���x"���,�]�<�BcQ�P�nЈ�"R�	cT����M�<YDc�r��1��Y�����F�<Q�ձP�҅����*
8�P{6�B�<鲆
(z8���J�%~A�C�N_�<1�!+��|�p!O!gƖkB�F�<��o	�;��B��[;Q�xYq��~�<�և�+}xe薋���b��d�Qf�<�!��.0� �a�=5l���
d�<��"Ι%yMX$(��^W$���|�<I$l[?E~*�l�!Ha�T�C�y4xF~8i�bL�qȂp���y�)�	{O�|���
�txf���J�ym �}Y�*#*��7\�@V$C7�y�M+,:Ѐ�JB�9�0C�gN�y(�q�:�$�M⧄VG!�T'!w���3�X,B���]!�LJ�.h�wD	�6�a�P��(v(!�D4 ���H�o"ʁY��ѻt�!�$!W[V��1΀! 1��F_Z�!��T�Ms�@�/��j���wFòk�!��D��(��&o��B�/E�!��q�%��O�2�&yz�΅�k�!�D��6��<	o�R�(�`�M�<!�ĜRq���Wc&V��K�-<!��yy�����b$�Њ�t/!��H�fؠ���0�����V9!�C�p}܈r�j��Se<���Α�B䉭W����KD��	 �3|pC�"Oh�q[�	 �j�h]j5�փO-�C�I�"�� �S������0��C䉴([4��BH
C��]�2���1˨C�I�3��c0�N�j��q��&����C�ɸ���[2��1-�Q&�̧:�bB�I.t*�]�7+W(8C�[�/Р"�2B�I�r�@�D ���H2���
B�UCL�⋀2:*�b�;|�C�IRU@��m�	8���k��M�BB�	/���ck�u���"D��!:�C�	8W%����o c~�E�D�î�C��
=�x�0�E��-"0�ˆ��7D�fB�	�+���ħ�bm�V�D�y�hB�I;=���+� >�@�1/�4+%XB�	�~0��ԧ�3[i.i�0(��sxB�I,\ ���d�ѵ3!b���S�BB��9�0H��� C'��Bh��)�C�I\���ao� �Ď���C�	;A�d5`���/}����C�(%�C�ɯmh|dZpe��o��0��-�eA�C�	��f����N�h�\�'F�B��C�ɣ;���{LG�s�r�
fσ�l(hB�I�v!��đ$8)F��� �Ju8B�ɣ�dX�g$�6%"��P�S�&Z�C�	��PE�e3}�]�g"ݯ~��C�I>�a��"�1zr6���"X3ZB�I!^0���"#�-<����DX�L�B䉛jwL��JݳM]�X%��`8nC�)� RL�6g\�F�
��f�%Z�"OmQ�2����w	I.80��"O����,���"��c�N�3"O�U��M�B��L�sȞ�M_r���"O��V�>n�A�l&X]+q"Ox In�>�j���	��v�lA@"O��Ct��C�����4E�f�+E"O��1�ED/Cb4�����`)1�"O(� ��bR�@��0���1"O��1BոL�|<"<H�Hq� "O�k��&S<EQ��-���%"O� AqВZ�RP�%����S�"O���cLa6���\Ȉc"OJ0� &Q�z��@I��[�_|��"O��V���:C�t��GB�U�p�i�"Oͨ�k�7���s'��1�U[a"Ov�+v-N3�j@��e�[ߚl� "OZ�b/2�tC1�M�dȞE�r"O8��O�#3�)YE�R5`|�e"Op�ʖA���8�f	�}���"OB�xT�L�P�a��7�%!�"O�8ش��)��t��닦,c�}�3"O�)��M͜�� ��JկZ]�3"O(���	�*�\XtI�xJx��s"O�Y[&�K�AT%���E����"O�-��-Q0 ���K@Kۨ\{XS�"ON9�F�'Tࢯʿ;Q$��"O|Uc؋e$�r� � V��}��"OHp�)��.�a�
�%O�� "OH���DG
�B4�q�L?D�<�*�"OJ���
.q�u
�9�>�s"O�K�%\,NHw	ή8����"O6�˗�SfT����/
��h��"OR5�A,!L2��OS1s��3D"O>q�&I�D2��bNح)���%"O��F��1&ʄ�#��t�#q"OX�����IZP�����3�X��"O^�U��ZrΔ��D���"OL�auGH�|�P+�Ů���"O
���Z3R����鑘b%Ъ�"O���*��? �	�hcܬ��"O�{U�;ø$�ceH�e.���"O�)��ٵj�����Q3'V�@�6"O��Ң$B�O��X�j�ܑ�S"O�Ds���4��R�hN�C��D�G"O��U�O
.1���SD�2��"O�$�R�?OH$q6/ҹ~0H0��"O"�SGF\=RY�#�A&�;�"O,hRe��9Lv�]�%�������"O\�s�M�W��	1��)�BP:'"O
y��D��-$�S�0e��Xxc"O��"�'I�pZ~=2�N�:�6(�e"O�1�7Y�i�PO��85����"O�)��͂&�ikw͕9#�2	�r"O���@�R�������'�,�i�"O8ɱa�٣g��U(sA@�t��e��"O2��SƐ(/9�]ЕG��I� 4�"O ��5������&K�h��\�v"OdiD��"y:�3�>*�"O\�K1�H�]
���
:<�P �"O��X��3�f!CvkFq�d[�"OD������RA^��ֈ$�"O������B���sf�G䨚�"O���Q�Y�8�
�{`�϶X1��ڀ"O� <�G�S/N��0��3M�,�R"O�T%*��x�V!z���|��"O�$r�)��=�l�j���
0�2L�A"O8���I�hV��  ���0�.�c"OT9rn��.�{h��e����"Oe�&o�$t*8Y1�9b��"�"Ot���6���b���bVb�XG*Of���̌����h�H��m����'9:ٚ���-�T� ���P���'�hiC�����K�^0�	 �'�>�bH��^�։8`���R�v=��'��5C���t� �:�ڶi�'��@feC,Sf�P���6F� ԋ�'�t�jb凌0��=Yu��Ky��
�'�pB����<4�$	�,O�Y �'P��c�a�7u�,��ۋ
!F��'Z.@3拌5gf%xg/ܟ h1��'�}y�)Z�=$!r�E�A�4�p�'��xx��o�& ���(w���0	�'ђ]yA`�)"N��"���Z�Ν
�'Q�������!��O�_�* ��'����a&N�{���ѷBR�<�'�@�0�c��,#PQ�4,̋L�x=�'�(J ̊�.�@[�`��~X�`	�'�d=`2��R	�mkƃ��w�+�'��� 針ϊ��1�OOTC�'�6�pED[�.�bp�ƌ�X2]�
�'� Yi�%;
*��E�/_k���'�hu�Ǭ	!f��,��a�G��\�
�'Z�T��x���U��͉�'H��#����xИ$�U_	L� �'�z J�*�&j7�ˤ@�6W��;	�' 
u�E��& ����"Ҍ]	z-��'TDQ{�!��_ H��9b�8�'�Xbc	4qw����!�Ϩ��'� �CmK�o�`��g����A��'��)(Eg?z��-�!˻5��mQ�'�<��Gˋ�[�H`��З7'�t�	�'��Hr��33Z�J�a�>#���P
�'@|	H�i2yN�@b@��1�	
�'�B��e�{�vlx������'�a�v!�+�Is�̝�Y
�'��djG� }��Y��K��3�'�v)�!i� 0��́r��$t��	�'L2���B��(�`'� � �"�'ir@�*M<nh��+Q��F` �'�nL�A')���ĉH?����'�d�`�"˘?+�� �h��<���
�'��q0��Ǣ\f���7���3Ϭ`�
�'�f�[���(U��`����#�$[
�'(̪�E�.\ԡ�1
L���j�'~E�s(*�ԋ���O�f���'��yp N�%f�ơ8$�ͧo�`"�'�49�i_���E䋘�8)����']�u{�l� �*�ɠ�3>1��'c4 v��@�T�JC�:�X�B�'� ��K�/��)�s�*9�\�	�'�$�
E`��1�tAYC��(t�	�'�0�j�D#H�<�ӌ/)��tY	�'4�C,O�=�<�g+׊5/���'4)ˁ��,։H��5�`���'X�4���X
G���iB*�o����'>��r�֊.���u����5!�'�A�(ON����NJˤ�+��� ��H��"4	�	۸rb��t"O9iE^�U<Mp֯ϲ=��� `"O�\�v ��0��E�3��\�"80�"OVI�
[�8p6MYG*�<X���"O�a#�+�o�H���F��Q"O+M��l4́1fO��{��W��!���:B���H�"A�ls��ޮ�!��T��*1�	D(y�(e�!���7 ������ß"c(���ʝ�;�L|�Z�����	�U���A0f��M���z�AS5}߈C�ɨ_��y��$��諤�;GO�B�I`�l�s@�"i��C��B�Ɉc]NL	�Y<,p>��B͍!_ B�I�"(����;�J�*ׯʈt��C�I�'q0҇KL�k�Dl�%���7%�C�ɘa6x(f-T��!I�R�JTB�	�no����N<J_ar�D��$)�C�I�~��D��A�$9X�H�3:�(C䉛62l�����:Qs���2A]t8C��
�QČ�uH�m�����4C�ɰ4,�9��/�}�DS��8HC�I:s*�$sB��}��M��	۬<XB��	) l�
�ϗ <TԽʁ�ܝ�\C�ɰw�,02��"M�dq-�#qC�I%A�4��2��=���a��U�[l2C�	kS�"ң?D�9�%�&V�C��#W�
e�aS=)R`�	`�`,(C��
����c�@9H7�1��+�L��B�	�7�V4��KD%���₢͇*��B��pT\���7bJIR5Ν,U��B�ɃG��8�3�WvP�ȳǫ�u�ZC��C�va�pIW6IfX�Y��G���B�ɯ�
���N�:J2&Ѐo�r\�B�I�Y�d����<#d��$�8D�\C䉾7ܴLRG�§:MrӧN�q)^C�I�>e �b,ؘld���a9U�B�I1>�,��<��T�eFL��~B�	��ؘd��l����i˅�xB�ɯwc``BƊ�9j�p�� ��>��C�2do�X�B���d4�u�˙nK*B��#Q��E�E�V�A)<*��\�g�(B䉁R��� iؿ6�+fě4B�B�$\�� ���҃B����M3�C�	L�f�2v!˙{+*����6{&�C��'^������U>Č:a�ȵ{
�C�ɹy`Jpɒ��	d׆��0��2x�C�2w@v�CƬ�-�\�+�f��D��C�0b��a��ϑ4���`�	y/�C��h��b�A9`���;ׂ_&"�LB�ɖ`���p��^33<xu㥍><�&B�	��Eb�J.z�H��h	�y��C�)2�H��L�Go�Q��JC
M�C��<C����E��N ���l��C�	�\<N��#�G�9�n�!���[��C��2w@L\9p'�!&n:�t@�t�C�ɸ�0���H� �5�h ��"O�1i��$a1�%��N#���w"O��။�=�;�N�dnI��"O4��1cM�{jY;��@�~4�[�"O����+U2�>Ds�,1�(�D"O�,��d,
� �LU�e�h��"Or�X7��'�Th�����Ф�e"O��
��ݫ*|�!�*_�{p��"OV���mځ-(Ah���fĭ9�"O� ��Au��!pe�r�#VmC�m�"O��B&D��qQd#)�졐P"O>�&���T�
	�b^t��E	�"O�������l��YG�&���"Ovѓ1IZ�~�B���<���"Or\�Ԉ��Q8��Ǌ!;�"�Ѓ"OL��"A��^�|���}�̴��"O�(��*ٵ5Ȳ]���="1�5"O���#Ip�Q2��E�1�"O�Yk�d��CtCƣ�tzd"O�B���:�d��vǏ��~�"O^�h��!�0�r�EQA�|ZT"O�e�b�Z�E�X�7ś�0�v�;�"O���קÇ ���c4��3	nd�H2"OA���D:]�:�+�dC�WevВ�"O��鐀љS�&�1vAD�j>pd�w"O�Ѱ7O����V�X#���%"O�|�$j�{[`��$��K�80�'"O��c4&ǆuw��'B� j����"ON=�/B�H�ോb� M�1[g"Or�
e���ޕzf���5�
ŨT"O���g ���}�a��6���[�"OB�Z>]����ɋo&lA5"O��2�.ɥ"��E�'��8&�H"O
�O�!|1�$���5W�8S�"O���皅t��p!	K�����"O�(���L}����+D��}h�"Oj`"��
�4YR�VO�"J��"OF]�f'J�~{���Q��-j��"O �#$jJ�& �1t,D�o_��(�"O�$��Z� �:�+��$<:�S"O��Z��7"M �2�X����"O�0rfhR;j��T FfE,�� pt"O<Ձq�٣<a��Җe��|��)8�"O�Q`i��~�˳N�M��E��"O�X��]!j�z�ʲg�$���"O�RQ���:x@�&旯Mΐ�%"Oh83���u���@��1r�b�+�"OBU�&e	�Wr�c5��rߊ%�d"O�[V%�	�00���NΞQ�"O�Ѳ3o[a�D��?mZ�*f"O$�V��/?j�A5BO�gNr�a�"O�Uk�e�xz��O�6C�I#�"O�����״��狊�ba)�q"O�����r8�r��5X����"O����Ώ�*dX�RIƀ@T��`1"O@R�+cq~Sw�֨_>�i�"O�ɘ D	T@��� ̯Tŀ�		�'�J8�Fo_;iQ��HS
�b9�'A*���+�
Z*�S� ��>�+�'�:�u�
~j���rg��	ޤ�'�"�b��$KU,t@��M3���'��8�H��dK��Q1�^~
@��'�hh��Ȃ���yc�ȶ�nL��'�(���8�ԅkU��x���K�'�P8��
LAk���.��h��`!�'��j��^+q����dgN^�4�8�'`�A���{��e񠝉P��h�'=b����b��%
Q�]�LRFD��'���Z&�@G(TK���G� �
�'�|�����<�8� #�P�r���'���5� [�p�oQ
	?Ҩ��'��iD�������E��t��'���hAe�0{A�]�@!��s�"O� ��it�̮w�X#��U�i���p'"O<���F]�h�H����E�)�
#�"O�H2�� &�~ŃW%I�i��8��"Oּ�Q~AZ��A]��M{�"O2`����;�e���<?v&��"Oq@
,0�H���9���r#"Op���h�R��%͜A�X�4"O�bdm��.�n :��¥w|N	sa"Oȅ����~8ȡA1��q�A��"O��S�R�@Ъ�����! X��I�"O�u� �0f�Z=�ꗆe�
pb"O���G&ɶc;���J��t��<��"O�Q�ggd\��(ң=�zm�"OL1���>V���Є�D�bΦpa"O�lS�m��?����W�`�
��"OPy��7	r,P���"�xʆ"O`�������X�=��Y��"OT�ڥ"�*\xi�� g{�,+c"OP�Pq�C�F.6�Z'��^���i'"O�����<O��Ex&�Z�Cy(U˅"O������z��鳒�!<O`�Q"ON���O'Fp����Ȥ[6�-XP"OJ0ˁb�>(��ظE)��T��U��"O�Ȁ�+��*�*%ZI��w���R"O�	
���R��D������c�"O���!ڸ��q*�ǋ�`����"O�䂐�@z�܌���K#����"O0��"��(Ј�j0-º� T"Obh�r�.+�0C����,E�̹q"O�S���|ء�&�$=�}X "O��R�?��[a`��/:� �"O<�;� �=��4�q�_�&��"O�XǤT�t�\A9E�ǒy�혰"O���N� /�0IA%G�u�Yv"O*c�&�t���r�B�T	� �"Oe��!�$9t��f�_�"�|���"OR`rv#LHH�I�i�4B�pLQu"Oڽ���� ^��E	�~�p��"O��AG
�>�>d��g��� �"OB����[�P��d� fU �=�"ONI,,��"Q�**a�*[�!�d�7:�d�V�Q�~�6����T�D�!�Z�A�ܵ��m�	E�bO��!�d��l2��#+�2 :�`��� �!���46(���J&P�y����	W�!��P�o�vMZ�B�|��1���!�C>^�X���{��=��얖o�!�ă�<ۼ�2f���I0=�JD�e!���(A�^� 2�Z�F�l�K��A��!��;wA�\�ש,H�� b�@5!�ϓ(����m�09�P`˽q!�D@�Gl���]�O��`g�1m�!���r5a%+°L{��1�Ơz�!�D
�;@X���N,�[���Q!�$O��$����b�ڠGX�,a!�f� ��X�~_�mA&@�$!�D���l5�#�JW���q���>!��/zV��I��mSԂլ��u!��^�rh����=q��sDMZ�Z�!��5Rz"@�����6DJ�Z
&�!�Ԅ8j  �d'�4D���F�!�$];��!4M�p���Sc�V$G�!����5A&O�R)>=q0$�!�d�6tF�cB�;r�Yc��j!�� �$c D�u�ʌ@�R�5/f�s"ObP�����C"��:P���*�0�`�"O�9�J��:�H�;��&U�
5�P"O���^XI�����9��"O��X&�֕F]�Dm��`=�"O�ŲEK�6=a~ɲ���!J�{�"O4\ɒ��-+V!��%g�#"O�%c�Òr di�Hج<|��"O�� �鄌uܘ�'��O�|�"O�t�/�R<p8���9�@��"O��QV�D�*>�h���"����"O�|Cq
�1�t��$i	(P�zM�2"O��Ы��)�q�Gǉ�SbF��"OB���  �   \   Ĵ���	��Z�v�G�4P��(3��H��R�
O�ظ2a$?�K&����4`��b�wa��2�� l�B��"#^
�7��Ԧ={�4C�2���:�'��&��(� ��8 �� �L6xT��B��v�`Od��� 0�O��_=	`�@�NC�^�p��Fꋈ	�,ё�\Cy®A�����tgI�����)\j�)�6�����W�8=F�k�΀*d�`g�,}�z1s���<��$។A�T)O`��D�ֆ ��T�ˬS���3Ҫ]!x3��� �x2��w�b�����$��'j���'�n�"�<bΪ!��EBdiBL��P��r�O-P�Q�(��|b�ҦL�x�@�Ѳ.�`�����yOOX�'f�FxB�7� \�%BQV4�p��7��#<��-�a�"� �,i���6H"rlH]��d�O�mh��?�'+���f^.D���������Rݴk^,#<	u-4�j�P���mU�}�ƜJW��Yg��q�Q�F��#<��h!?� �`�J՚��>\�����`�Gy�dVD�'Z�0�?�R-��	�sݏ���Ќ�Qլ#<�0J%-��d}50!X��[��3�ߌ�1O�#��D�!��Y��т&����h�@�>
��@��6Ŋ#<y�F'�I��
^9���;� JDb�S��'���ӯO"�y"�(_�1�|aa���y�×�#z��0c��;*���Dj����/P��r�|⍗> �@J<Q�*.rcJ%
�G �?H��MW�3���rTf�e�	h1r�C��4�Ie꼼��U9%��Řu�Ȝ�c��XB��;��  �$��U�<��C>A�qt�V5��|hG�g�<�@cE�0a��+z�8w+�K�<qTaU�D��p�lФ_z�����G�<a�'־P�b-�T�P>�(�@�G�<a 
(@͒�z .��?
��1�j�n�<��&=lH i�bI9B�!���n�<Ir�ƛ4�̈@���!p�!@i�<���Ÿi]L�#J�P}�����b�<IRB��"�!��	�Ĩ�wD�^�<���8p 4�J�u�N�Cv��Z�<� E�d�Ҏ��!`�� y��RT"O�p[ŧ�޼A�4�@m�^\��"OX��H �2!z�� � z@dxҔ"OF$�U�ܳ3�D���h�7|�jp"O�;� \\�01�G�	���9"O�	)����,-�p����R��A"O���f$�>Bx�)���	��"O�   �  o  �  �  f%  .  K4  �:  �@  G  WM  �S  �Y  `  _f  �l  �r  (y  i  ��  ��  3�  v�  ��  ��  x�  �  �  �  ��  +�  ��  ��  4�  (�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;����i`9"�ˁl�$@��- G��D��O��2�	!0L�Qd�*��PZg"OJ�R������qE����Li�"O@ӥg$x�|���ֱE{�Q�"O��"W����i��ۇI<���"O4)遪@7��P�����z:�!Y"O6�#�`��U�|����%(@"O��J�΅-����		���	շi�hC�I�(���Q7n׭A)�� ���G22B�	�{n@ 8%�@��j�;(��!@�C�	�/���#�"[���@(K�c�E{��� &a����k)�
Da��>�~���"O����<A)
H�B�%`��i�w"O̕(K*$r�"�d̩�XС�"O� �fn�-V�&�
C$M&0��RT"O���T�'7_�����߇ke:%��"O\6�&un���'��V��
��6D��xr�@�I�H�j�O
<��x��"4�	}���Oi�s��Ki����Q�7
XJ�'��|A���{JT���5�
�b�'^d	�u�Y<��k��}e>e[
�'*j�� ��,3`��{�[u�m�ش�Px�E7Q�I�T�[�\���)ȫ��=���|�!�-%Z�xf�@�N��P�d���y�E�0P�ܐ��K(L���;R����'cў�Oz4�c�Z>��H
�B�Pu����'���e	ݬG�.� ��>P���'� ؐe
T	v� p��_�R;�'��<��ǔ&�v*�)T�AL���#��;"� JC@�X��L9,0�@��"O�u��"FKT�D� �ԧ}�h$""O�h"'�;Hs�Sdd��op���'Vў"~��&L(
m��nS;#g���¡X��y�W�z�B)�֡ڞ$�.�������yH�jT��ߑ1�%R���0�yFR�5X��]�$��,���y�)�6{���Fj\9N9bT���X6�yb��@f�\�Z�RC�߀�y"��KN<�P�O��+J� ����0<Q����)+TX�i�)�d7�����Q�]�!�E�8���P�	�<F٢6쓃$֢=E��'-����@,S�b��7��`H$z�'���/�r� #TfΞfE8yK��?	� ��3��.BD3v�/�>����H�MY�قG�1c?zib�e�8ʒB�$q�zA�''�m�L�?J�|��O�"~J���/�  �@�ӫ�"J�I^I�<	e�)�8D�A���MM\�	PdC�'��yr,G������C&�Zr�E��y2]%B�F��S.˚<�`�Z⡐�y�����������"1��أQ� >�O	�'NQ>9�0װk��18�)+u~mɧ!$D�����p#ȰR(�<=ެ��Se�hO�Sb�)�Ma�
R	��Ԡ�LK2�U��nNZxB��nՖ` ��5�hd��O*]
R�Ӵ �ia�F�GbJq���D���,i�i��9+��PC����!�M1Yl�)rfA�L�L=�H]�!��	4��a��,ۊ_C�ecwf�<{o!��B��j�S�ȧf#�p�$F݌5X�^�h�<E��4O���"$%U8���Ýzsb��ȓ]�~�bh��J��1�SZ��}�ȓ
V���`ǔ1J	9e�O.�8e��I�
�v�R��Tي@M҄�����ޔ�y��=R1��Q�>�<$��8�y�n�e�Js�"G��h 1aU"�y�d���Y��)9&�]��2�y��� ��U$�.;�虹#A��yˇK7`˱��_�p����yRF�&s�L�X���N��y�6eǍ�yD��{˒��F��� z|:����y"A�;p!��`�VΌ���'�۰<���̵~����A3?��!
�����!�Dә~�X���L�.�xIyVQ�c�!��\���8ׁ �<�.D�C˅�z!�� �B���ndt� "G�T�tR�"O�LB &t��]ZP P/O#N[�"OA�Gx�����l��I,�a��"Ol�����-! �@��I&3t���"Oz��e�(o�2E��gH��1�"O5�1�+>ꂬ��L��_�e��"O`��5��#J�)�3��(�֩�"O�=�s!�c^t� S)�q�Dɂ"O����v�n�Kc�������"O1:3���,8�u�@�S1�ّ�"O�xjW���4�<��1ę
*����'���8���\y��`,A�i� h��3D���i1)��K׋Jd��TR"G/�nӺ#<�}�PB�d��Ђ҅�F��a]@�<��k`����q�]x�t����Q�'��yrj9
�ہ�ĕI��ڥ%�(�yں�v]+P�J vM�8����y¨�Q���
�>k_ ����ybD٬Z���@gG1cpuZ�ɔ�y�m����J��@6k�`:'˟)�y򣀿��U�F�ZmyrP�L��yBf��=~���cV-c�4-�F�&�y"�m�11p �)^[.�ň϶�y��K/�9Jpd�JЬ��)��yB./M��}���2F���# ��y-�*�	��7�������y���8E�Er3���'����D��yB��k�<��w�"��ӬC4�y"��/7X�RD�j�J-�r��y�7U��)&̒?s��2L^-�yR�H��U���X�W�$�h#S��yR"�D6�E�&~��E���y�L��14��2咿"7D���
�7�y"GE�� �#��.J�Q�K��yrN�9Y��:ebR���U8!��yRE�]�}Y�!~J� :����yr��=	NI�u�D�!�8ʗ��4�yHI6�zb!�	���Y ��7�yR��r�V�����
>��H���y2��" ��ܒ��ԛ"p�����yR�
!J�f�Y��	�\IҊ�0�y���f��2L�
㔍k��A��y�F�:sx��+�����siC �yҊؑ��M�2�� r�X �m�yb�5a�e���X�.��*��y���q�| :�腼9ْ� ��yBEϺI��Ȉ&�֗8<�@�F<�y���(H#�X�z?(�zP�Z�y��(E�0%V�K�C.�21ې�yb�D�Q&�۷��8J&u���)�y�x�X��膛9����
�ybE�f���%�h΀����y�k?i�̺Qώ>=������yR/
g��@z�c�!e�(�]1� B��.O������tm��җ+"RB�I�~5�wHP�Y ��V�V�NUB�ɁRRͻ׆�"*�T&¿U�C�ɳ(��LPU�S��Y�_J��C�	�tx�QB̗A��c3bX/)��C�I*aC�]��Fߒs��5Hv}FB䉀5�����i~k�ꔟqQjB��K%{�`�>m墵�B`_(/ݤB���A`�.O��F�
���3�xB�I%�!+��X�Fi<���Έ,,$(C�)� J�c�O;}n-�$�N8E��i!"O��z@��t�N'@K�h��q ""O�*3쓳1�	�C)�2�@�9�"O6tA�͕�)�A�'>�=��"O �0"�Mb�%��8[y���'%�'���'$��'e��'s��')ґ��  Tz��# ��vX�4'�'��'���'w��'e��'^��'*���)߁9]N�����<V�QW�'���'���'o��'c��'"�'�|�Y�Η0{���6
��j � ��'���e�i%��'�R�'���'f��?t�X�(s,N9j2S�@���'���'��'b�'���'�b�'݀<
�^�Aڰ����Ɓt�"�b��'cr�'CB�'�b�'���'�2�'m�4��lX��̴,��(�K�7�"�'��'���'���'�R�'���-��� �ϕ)��t������'?��'���'�B�'���'�RMY����)�.P��<i��>=�b�'`��'>��'���'F�'��J E+*0�d#Ӯm������E�B�'+b�'�R�'1�'{"�'����4NyÄ�@5�d���X�)�'��'O��'tb�'�'#�g�43l��&�"b�2���VP��'v��'xr�')��' r�'Z"��&xܥ�̃�kV|u�M�Xr�'��'��'��'�T6��O���XT����,X�b�jq�#�öy��q�'@�Y�b>���&�G,��t�N��K����a�*A2z���Oz-oD��|��?Ac@T/T,�«7?G��s���?���~^��ܴ��$v>�������/O������R7F��`��� D b����fy�퓜er8�ʖ(H5΀Q�m��/g��ܴF�&M�<�����h��Κ� �\ܳW��+2g�Y{���r�,���O �	u}���$��b��f1O0�;wF�/����$�%Z�����<Ox扽�?�U-/��|��)���8���A3�E��F�sC����d*��֦͚�l"�!n'&��7��~���"�%f��?Y5R����۟�͓��D�6K�PXQG��A����;���xI��v�c>yA��'�����e}rӒ�	��n\�r#�)G�l-�'����"~�*�f��$���p��iu���Bg����4��x�'h�7�-�i>�!����������5j�q�����|�I�h��en�Z~25���ӀRg�9�-��e�'� UP�y�'�8�a�eB�(� �K��\I�n�r�'�9�gF�o]�\Z��D�h����L@�Upz(y�d�<bti�_9k�,t9�%��}x���A�|��E�GOG�I
��B�#�/JJv� ���}�Y�b��1~JZ(�g�(Uy8���&brM�f&�9f��a����i�H���?bYf��U�ĉ�R�#$�8R�N Ǣ�b��p��ʧ�0>�FF.rx!!�ω�N��}Za��v�<i���".��b�K�*z&��tl�p�R�c��,��`���A�Б���#3
�aZ�N� Rv<��o� iz��ӻLM��s�E�Rx$)��mj�#1����$��N�6�:b�ح`"Გ	�Q��A�톢5����	��Z�R���麰k���{	lXS㫅p���Cg��-l8ېn��|L�����2D���q�� 䜝��������C�	"wTLڇG��\i�}�烏7Z�B�	2U�-#T�
�(�1#�'&T�B䉷Q>�0���óU|��{�(��pE�B�	�G�����1l� �Kܔ!#�C�I�x�h�E.���A`$hբ�`C��2}��)�+P-O�P��1O,n�dC䉻SXj����'�qb�ΫN��B䉣'-:��b
���l�-֦B�ɲN;��$(C،�FN8}�B� NI����"��iO��DB�	>O�ꉙ&�_�=d�H�B�nv.B䉼�L5� Oއ&�ݘS�U7m�C���hE�s��4��4[pH	�C�	"` t�JG%[=
��(�&�-<C䉎6�b����H��s6͕5H� C�I!]�2����Q.�Sb�֓2RB�	��l��ȗ/4�	�֚��C�B5d}�(�7]3h	;���&D�C��	a�\ڱm½[r ֈ�Y)�B�	�Yˊ��A�u	˷�F�A`�B�ɚ[��U�N��c=Q��ȅ�C�	,��l؅�ɣR�4� @E���B�ɾ^Qf��S��&|�85�!� f�B�)� �0c4�Д�f���iL'	��y��"O�B��G� &��Jo�����"O��SV��nN�"��o=z5��"O�e+��՛ ���"C�ҝ 7R=�
�'�j9Эځ�0�w��YBpi�'���c�����$$5	0�Q�'��c��p��2IF�6����'N�t� �
#g��9���	2���
��m��u�4�ТU;�a��G�{�h�rg�S��d���!��e�|�*b'��|7�>�VrqZ|RB���b��(�O�rXaӮ�;m�F�i��%c �	�'p���1?MX�$E�Uz�u�'-����P�e�ReZ�OI7 �"r�C���,��Mָ~�|Њ���n�<Q�eD�s�B@a�DĖq�*�h��M	u�F;�'f�Dm�R��ܕ��O��H�0t�b��W��_��� @�'�J"A� =��iC��W�jX'LԀ9���h�+[�v�*sѡ���0>��FE�5��\�E�ߡk�tp���I_�'��Slz`�s�� ]�r�{�?���8��W�i:�s4؁yq"O��8uGY�V�c`E�}��ƾi'�)�˚� ��铤�Б=Q��q�t��5�!�$����4LV 6������ͩ�y�&2��M�d��Y�25��O�!��`#��lӘmq2F�F��h7\?M��:p0Ġ�����5�Ã�a~��Q+�Ԁ�Ղ�.5t�����+�����AZ�Y���PG�{����IE��EC�+U7��87�D�*#>	��Ù(�|�(�NͱYgF�r�P?q��/X�؝���4JzXh�&&D����"w%�(�&D���ti$Ji�,pS��/�4�B��Y�"��	���O�e6���(����3g$G$;N!�d��� �( *�sNx��ϲ>�&�����e:g��B/0�[ҏ,Fx�f�5"iT��e� \ۄH��B?�0?�T���ws��0��.���D��,}����ɬLs<��%H
�Ta}"��5>z���ɔTt�2C.�)ֈOD����W/1B<����=��d�Oܖ�H�a��~1Ն߇����'�rD+	&K
j9�s�^
u1�xڜ'4�a�����~G�RK��7�?1�#�Q	@��l��O�<���)0D�$�V���rP�@�bX��3"$�<�e̫!�2�	3Ƙ��0<�&���v�lK ��\��q� �pX���	% YD�Ҧ�ũ#N��84*�	Y��
���-_^��#��#��\~��u�6���)$�LDz�nR�Q��X��)�P��kpX4 8z�b�A�/!!�D�6��h���4#Z�#Ʈݯ	���M>v�9�=E�ܴWz��	�0sp�x����4��I�ȓ	�TI#g��\o`9�������'���x�'6��Q���Fς*6�B�q�춄��6OT��u�W�8��dQc�.=���"Or����/D�4!�΃&N)#��	�-���ق��*�:]����-m�r�k���=�B�I�jm.h��˺? ���M��6��%M3�a[���s�
cd�"�:EŻgD:���"O���@8HQ�)�LI�Y��_���D�
��e��ɝG��|ᒆ\�d]| �� #�$���� c $�{�|�ܕ�#��� �$��Q����B�	�V��a�� ^�D��pQg�R�V��'	���N�L`�AF���6�(� 1\q�� �j�Ӣ"O�ib��]F}�pTb�2��]�0�'o��R��J �??�Ϙ'��i���u�,�1�Ewd�0H�'4�k�GW�v��hP :nZ.|�rDT	%�t�4\�]���''�I���3s�jq�#� 3b��	�-E���R����uj�$I�V�b-L�!�4���ڒ\C�L+�'��0Up\ɲa�ffVQ"�O๐a�Ty�f �lo��D��c�0q� ܀��� ��i
���+�ymE:g{@��K�C0�u�vBC�����=�r����S���~�<Q��-0��;���"��L��) ^<Q�ˍF �0���#1��Qc���V²�oZyy��
�\��N���DQ=	ANa��\m �ej0.�axrS�/v�nԑ� Hp�L���d#'��U��B �i����	#�O�p�GQ�z̪G_{J$d����Q'����3|
�E¬O�+�L�?m�tM�^�u��fȨA��V�*D��$��M+PE��8���!Jh��۰
E�j����d��?�Q������Q:`�ᝡ[W��yf��[U�R����J���&7��ř�hq閼i���I{���:7�
n]�4��'q�n#<i!�2OW��S`'N�}��$�s�'&�x��e�"�M���r81i%�'/vQ�s�ʵx0 ��j�D�\t��j�}�]9�p������9Hq�AOAa�>�D��/R@�!nZ1TV����������<ͧpE����0����� �(\!��$�\�3�CD�@)9@�3'��@F�3�D��X�p�s8O��e���{���y7I-R���Q%BC[�����!���?a6g�$�58 �X�ZH�!�ɢ^v��fM�C���Y��c�V��S�H��#<�3���MH��� ;{��!R��D�'Ul@�$w��y���/�I@�~S��*viعzT��y�CKc&TE�3m�̦9S�Zt� I�cز\Y�����X8<&����ȧ>��L�-,D�dD����~��|��iA6;�J��r������P��K�<��b%S
� c�^������Q@5=O�t��IH~����y��W�p��:���,Nf�Y"�G����?���ˏ~a4�`�b:�����gSI��lB@G�)�~��'��84� "<�Q&��S*H��Y$�X�C�$�Z�'�t�PE*�56H"0
�"������h;l-�d�P�v�b2m�.]�	�m.��Dǃ��y��'S�s��а`�*m��I��B��%�Th��1��O��PĀ(�?�:`c��
�@�!�޴F7���#;0;��Ն
���Lip��<�����t���g��CEm՞b~\�jc�ߥD�B�h!�EB؟�J��ʊ}H
�[�σe�Q��8{I�����5��=Z�!�O��
Sj� 
���/����I��M��и<��"T��~ң�B;7��	�/ �Zy@	��M�<y #˾W����ə���;���q�;v��9p��쨟�hE�_�s�Y��S j����"OT8�
Q�q�<��Q�_K�m��C��������h��$��j��mK�ΆX�$a�� ��;�!�$�8R�;Y#�80f�¶)�"m ��`��1�'�VXڰX�5aJ\{$ W��Zۓ+�"�"1+�$� <�R��5�jl���VJ:!�$���x|�"�fX��*��ұO�H�-��|
��E��'��R��!�oػuV�t��j�ykP-y�0�F!�I��jX�41�������h��$^�Ԛ��f�Q�P���j��E�!�D  y�腡(U�� z`j�:4��	� )ҡ�
�>?B�	g`N;hGr� ��pӦ9�1M#t6O���F�
[3��c���FP�I�T"O6L+�KX�w��ع��6�H�J��I.��ɉ�鍮1��1{�cϐCP|� �*ӈK]!�B/AyˇNɼ� ����g��(X9Pb�"~n�2?�R��RF��py�	���72��C�ɻc*�K�h�R�L�"t,�^���{0�1a.-|O�Ԣqb�;:ԑ׆?Sۈx�7�'&��c���M��O�>HL
@i\�����vn�<�ä�4�&��"oI�qLnpJ���C�'o�bTD��H��� �H;��R�*�	eb��;U"O�H�fb�)v��\b	'J��p�i^��2�"�u�S��M�b��@^�,����T�L�h��x�<��`^��p��b�Z�Y��l�s}��W%k���ė�OI8<S��+@@�3wo�>h�a}b��v扞)b��
M�S�\<2��U�B�	�.�Bp�Z=_�p˧ �%+�#=YeU'�?��v�]5[u��`%�<��b�8D���:7����0���.9���w�@[��M�S��M{����&f�LȐ�Ӛ�4����n�<3�����%p�F�%CȂ�xƯ�k}�'��V����M�P6|}����}U���c,�dK�}b$�=�~��Y�d��G�Ҧ}��@2�y
� vq��rM*L�����Z��`�"O1���2T��(r�Z4f��Y��"O$p���E�6t�P�B-�l�#q"O��aW����]Ѥ�]2ZtF�aV"O.�`æ�(x�:h�,�fX9Ѥ"OPI�7
�!e�|���NHp���"O䝛ǭ�mT�;h�4[�8e��"O�,��јs��|Y�ś>ʸH`"O�Y�q��,[,�HG���tv"O�a����dal���D������"O��SH�;�~i@�f����'���R�XVh���gP�D��L��'Px��a�c0���g�/l�ER�'�>�J����tٙ�!�$���
�'G�=5/�9�eK�7
0k�']�=kd&3`�QEA�&e���'��:'D[-v���H.
t���'b`X�r�,<FX�ABړU8Z!��'����Q�N��I��h��_!pt�
�'XЈ�&�/%Ҋ�QHɯW( ���'�����e��I`c�JH�u��'��4���� u�Θ�d+K:	��'30�7'�).���^�1Q�}h�'�<��5�ӞB�"�x��-xR6"Oᓑș�r�kFڡ�i�"O��܍nix̉1�|`#a"O6-S&*ə0x`����?`�PI%"O qx���
e�	1��;W�EZ "Oڅ�׬�7W�����6U�%c�"O� R�7�@�B�n��،"O���n�6�4��-ۉ>�b�	r"O���I_�4��]�m� =�ڰٗ"O 
$!��*hj��H�S3V��"O�=�X���Z$Y���3"O�A��E�/��:((n�Zq"OT�@w���w�-p�X��bM>0X!��@6�P���-��՘c��+bI!��^�C�F���
�]��в	�!�d�3bК�S`bX43�$|��͊!�Ď= p��T���g��P����!��I����+pj�w�`EaLZ0g(!�GP����"R<fiT�K�(��&!����6��$Ό/��4a�>)�!�B/(O��k`�������!�_��P�h��Pd�t ��Ь/!�d��	e�M��-^�>S�8zvj�	�!��O3Ծ�����8FԀ��K�-	!�!��\��	֎>���H>M�!�Z({T��:��ˤ(� 2�A�!�dQ�o.���ݞ<=T���d���!��/i-�uP�˖)�Z(J��W�!��Bs^v��%/	+#��r��k�!���$툴�De�2#&��5j��r�!��& �}�3딓F����&�,�!��ڞRb�쑖�H(t�`����`!��+_�@��[�Fgd��CU�6�!���0�2`��a�8y閉1c !�$X�*��H�s�_�Pr�U�� �r!�d^]LPR%��x�b#�.��?�!�ė%)N:���%H:�|�U@� 5!򄃮o:Μ�@`�2G��~�\�'����O=&��&�I����'}�	��aU8C�@�xF�{��%��"O&U�����G�l*P,�#* �A"O� DMh�F�Z`i(���J�I�@"O�p%ʌl��M��F[��1"O$��-�*$�Z�h�)c?hux"Oh0*�@_�<�f��塎�6Re�#"O\��b�-{���Ч��G��Ћ5"O,�S��T<4\�y! ǻK�D��&"Oڅ� �T|@�/�#Y��l�u"O�KcV�ml�`�:/��4Z�"O��q�� �ƕ0��vyޔ�"O@#S�Ϩ�@)��>c=���"O�p(F��u>�IA���;|4�"O�xе"��+�0��ُ�Э��"O�}�5��J�NHxg▣a즜��"O"4�E�*Q�F��� ���	�"O�Aw�V�f�6�P�+�����"O��@&��9���@��b�(bF"O� ���Y�n�  ۨ=VJQ�!"O�y1�gT�cT�� �v>,��"O@9zƣ�aTP�����Œ7"O��V�S�x�z�BE��4��p�"OJ����b�N�'+�0�┚�"Oʄ�����b�t�gi
�z�nQS&"O��M���R��W���|�,P�"O�m�gn?|���B䇷l��p"O ����7��fC�0i�x(��"O�$2��֤kNܱ�� Kh�qkA"OZ��.�9혭�� N�]:c�"O29Q'�]�Xy�E�`5�"Oxd������$D����<}p\8"OؚU�-�{W䒎6|v���"O|@rw��!6��3CS�o����g"O�)���0\�ɨ�O�]ap"O,�z��ܦU��,��ȋ{�n���"OB�x��E3 Q��U����`"O��R�G.i������+0�5��"O�����/%#�x@���),<~���"O���t'�>!\ ��9a�ۗ"Or��V�E�����6/��"O�A���T"h�q#�6�%��"O�����E1#!^�7�fp"�"O��;���iQ�M`a�ղP@q"Oza�`�W��D˂�F�S�8�6"O�5#�6��4Hb'�=?D��"O����J�Z��Ʒp>�l@"OȅB4�ҍL"�I� ֝8�T�"Ol�%F�L�����nS� p� u"O��ҠL2v�<xJ0K��$<̳@"O�!��K-J/��b�)N P�r"O����d@���IxǇ�>' #"O�H"4iԚ.�0�2�fC�r��`�Q"OJ	c�ˏ����p�[-lԎ�h�"O*�S1�ŧL�~ �bؗ3��=C�"Ox1��O��_{.P���ڴt��ѻ"O,8�`�XP�C'�
�g���"OR͋�B�>x��!��4�f���'-���ԮS+ �p��4ɆQo�I�' �5p�G&+�4�d- }�tB�'� �jc�݁W,}�����x�lu3�'�@�&�#a�Լ9$f�wF2qZ�'�t���ہ ��Pc�ov�`���'���C̋*�2Xin�oPT\��'�xy�C,]6.�R)�qf�3?����'z�x:RL�7'�i�g(Ķ&'����'C.�r�B�tyw`�i��a��� BE��N��m^74˖��*O�5ӥ�ˇ[K���`خd\<̩�'�zႄ��<�h'�T'[e�mb�'��-zC�E�k�d8�VĘ�_Rk
�'o��R�^1G�6\�&��R��'M�@+uE��D���&�"p!
�' �)�M�7Z�d�X�h FŶ��'������=m�R5	�/r&���	�'�8��Ӯg�p�P�_�kJ2��
�' �=��A��va���éQ��dP�'�B��ٝM*�$2`B��(��'_"��d�ֿ#p�t�'�^��Yi�'pXqї��$N�`����V�@�'<���,�"\�rؓ ڐ-!�=��'4\<��g
�DɈ��)��OoD�P�'�$����\�K��M��:����'\\����O��=��$T��n��'ݒ�y����R���5@���!�'#N�j�n�O��@��,�rd��'�t�c�S�QD�A��L�V��P�'���@EO��Q��U`�K�x��
�'A��
B���B垭V] ��'ӆPZ2�}E�I�L��\="	�'�x���׬�by�en6����'���"���(I���'�Hi�	�'K�-�e��ra��
 @j��0	�'O����N�T��C��7@ eA�'.���tG�3.?y�딛�uS�'�*�A�A#y�)'��:~�"}��' �T��ܶ	`���^�*1.m�	�'S<�Q��'@n(���l@�5B�'�����L�#ˎͺ@L c՘<`�'���S�ʪ�,�{`	Y^in�8�'Nb���䛔L�@���n�2[�2�'I���+}C>�z0f�)kR�d��'�­,�=��i�" PX�<�'�� 	�M-}��	��^.5ʶu��'{��AS��,�LY Ύ7��t�'H�i«��z�V 1�x���'���˕ޗ6(��s�V&?fF�9�'���#Gʘ:�L�Ci2�\�H�'�Ґ�dh4zp��R�"U��I��'��Re��M�p!u��< :
�'�5S�E=V���C�	 �l]Y	�'��5�D�5_,p��ʓ�4)	�'i���� �G�8�X"+�:]Ĉ��'� TY��+f�v\�Q�^�N�D��'�YzVY_I��*���
}��u��'��C4-A�B�h�� �y�����'���۱M��.���RIP6�a1�'�d�Z#��?SH� ��U3�4dY�'ӊ���W`�<��1�N_����'%���@�P�H��8�ʍjR���'�hyxSo�}8���ޔo�8��'I�9C��V�M�4q#Ю2���'�l������GhJ��l�&�1��'5,���@�0�`�afFޕ[�� �'&�$�S��T�☀��S:)O`h!�'y�##�t���@F���W� �'1��b�-��%0A1㤆5W�̹��'�����o.%������6K�<��'���A������K�a�>C�����'|�Q��վI8�ae-Q�
�'��P*��L�B�ȯ&Xf���ô�y
� ��
�J�6O<<�A�30�qD"O�EK@KЊtn��Y6-H�X��\� "On���R�XDt*2L��(R�	0�"O�]�b�G�rEN	׫�>8���"O�x�B@�1o��P#�ѫr�"03�"On�'�#rpڅ�f�˿k���c4"O���F���:4��ɐ2�dq/�!���(x֌,p2
	obuxq�2X�!�ē.U��H�B��m(�ቄoS�B!��P9K�@��V�Q^z�Y$!�� �!��%g�uJ��K�`��,a2��!�DP3J� �*N
{�X�BnP1?�!�$�\�i��]�}�8�ycك`�!���Z9��)�<(�V�#F�[�!��ijzY�!�� �̈藠͌p!�$Ɲa� (���цu�`����מA'!�C4�y�2�߲!��A�r��-w!��S!}��$6 H��B,Rƍ�_!�ڬx��A�r@P�%w��y���F�!��A2`Y�C\WR<(ᩉ�_�!�L��yv�ěHr��v�!�����&�ϞkB4��2)>Q�!�d�"�����yR���.����'��jM� ��]9aC���@�c�'8�H��'Ҽn�"�sS��*}8xz�'�D�rSȝw��I��@�HiJ���'�Cgbճ&V�AJ�d�j��i!�'��i���7~��Ќ�?d��б�'#����>�	�$�ܴZ7YR�'�jL����Hj��g����'J�b"+K�S��!;�*ѿb�^��'*vaB�?Q�tbwѨ�F��
�'jᘰ�ƥhwh���-ƢW�t��'ƪ	��ՇOph�+g��$TL�1��';��Qo@�+�)����"�p��']�x�"kQ�t�2Mz����-�3�'�*\+���'��ؚ�d	r�40�'{28��"[,�[f)F ~�A
�'�4�aᇅ+�����h����'�l�q��V�P��SbM�(!��'�:@3Ƈ�C+ ��H��X�1��'�Y`�.\rh���.U�����'��T��LA
K:�r�M�d���'�"}� m��BP] $�I;pmY�'�$��nx����K�O���
�'��Y�gB�C�l8�c�:��
�'��C���rM����0�	�'W�ܨ0M'"|mH��� K���'\>e�W�O>:�X0� !q��[�'hЙsU ��@�*]�".U h�d���'�sw�va�염}c�a{�NP9�y��UL<�3�O
o�52G���y����?BhP�׬�gc���3�y�"=�(��Ja$��!DD1�yb;�Ht��0%p�\�A��6�y�ϋX���+u��R�L5Z�H��y҄�N���$��*K�-���Y�y"��<�NL��!:�)�v/W��yr�	Ln��̈́(:1Z&+�yb��$x� �@�6�����ͭ�y� �?|%(ŌI��M�#LL��y�Ç'V9��� >5��e���8�yb�I�nW�3�倒1�5�����yROO1;}��8BΝ�#��ٴjϛ�y
� ��1c�*E�L����(I'��$"ON�Qp'�` ���m�}08IJ�"O�*�H��/� 詆Ʉ.�%	�"Ol�8�A�<M�6��̊�>Jr�rA"OxA�N�"5>`U��k�e�lp�"O
P���:>�6eY�I@'U�8kd"O����y������` �u�"O�h�Ϣf��p�Dr�2-��"O�]ɡ���p3d��k�b �e"O�I�Q��1��Iwb0v���"O�y�J�!R� �A!CW�zeX��"O�p
��Їc�c���tN�(�4"O�58�E����ī
m/eK�"Oچ�ĕ!��E��#B&"��h"O>e��Q�Z�zQ�7���"O�)@'�w�81C���+���"O2�hgFX#���w��"�P���"O�9�T��`�N ���:;�
4iP"Obe�		dAr�@#'�U+p�#"ONX�(͚-�`	�L*-~�l!3"Ov�z§�R�vx�+L�v\*Xt"O�Q���r4�K�L �p���T"O���S������K��W��]�`"O��p�B�,<�b�ː���`��"O���C�O�$�k�ʖ�0%�ݪT"O����ڠxL�@�ƒ$H�=;!"O���l��%�Τ�Q�}��1��"On��玆*�d�Y%i��V�����"O�P�U
�VL(qHZ?>����a"O6a��B�c��܈�f��j,��"O� K��Y���j��8��Q""OF`��!�5:�� �]�'�B� "Om	��D4 8J�e � BiH��g"OzȔ��
�hC�O�d�`"O�U{��WJ�&=��-KZP��˷"OEhE٤?����g�ڃ"�� 3"O�u�r�N� %�eA$q�]��"O8g�ڨ
b�q���zb�9{!"O2�km0��Y��Z�ư��"OTkBl�"5et9+S퐃=�h��"O�ٻs� ���i�̏8����"O6�2��ڸ%}��+^��T�Y�<A�.J����&�$m�Ұ���PS�<����K�z2�Fzn��&�X�<A0�V
����N�����W�Y_�<�cu�8`�힀$��-�	�t�<0NT�sW��`�#ٗ7�(�t�Fp�<qv�^4I������^T�񣤉V�<ф�jCr�X3G�<'�xM)WS�<�u-݀,`l<s��6S��0#ʙO�<����̣r��>\*)�rD�<m� ���UA�?R&���aYK�<)����X:�L�AT��扙�OL�<�1'Ā��=�Q! 9%��m�A�@�<AS��	c$�x�/	 C�$dQc��V�<Y�A*6���@5�J�"����l�G�<�7 B23�|ȁ!��~'�]{��G�<!�Bi,�1	*��S�h�<�@I$t/H��S�·*�ԩ�nC|�<�.�54����E3q�����z�<�5g��|y�n�33zT�,Y_�<��e���$��� �?*\�7/[Z�<yQĞGJ��@���,<P4�"aC�V�<��I�+	g;�*P�x����7��T�<� 
�y�ĝ;t=r��0�X���q*T"OM÷C�J�*}�I��6r�}�u"O�M�WO�5�j@b�<Yad�"Oh���@D�BE+ШÔu:`��&"O(�Z)��C"cS�*"��&�y�<���E#���R�����)v�w�<AW�ڃ7V�j�����Yv�<�1�dq�IF&�~�Tц��G�<��@/06ݺ�d�m`�3�BY@�<�Fb�s @��D���
� �y�<����49΄�G>,�m�t�<��g�I�ƭs�(�t3����@�j�<�^� H��kgC�fe�4����d�<97���Uʨ�	1�BpBz0YQK�k�<�r��r�|i���=�0�ca��S�<�#�R����	;�Lġ�Ǎh�<��D6���ҔL[*��t�2�O�<�b"�6+xA2Q/'y<���a�<�A茾{�u:�K�3w�̀�h�<��i��|���(��D��(XC�A|�<i�e��:k�2�+ ���ţ�f�@�<A&�"l^�Q	vo��h�@�c��T�<�sϘ�a3�	�K��ui�����RI�<��eS�B�� �b�20<������<iR@�3d�p�p��B�)�|��Y~�<As!X��=���U:6��dK��TT�<ipf�5qJ�0êH3;frh�w/E�<����&���,M�iW&�hcJ�g�<����):�f}�$*�{�*æ�`�<)E��-~��3��A��.Ѫ�`^�<� �4���i$"F�D�W.\�<��Fsюt����#z΄�dD�Z�<��F%��P��� ��X�<�thN�jg�Ѐè�r��%3�!JZ�<����$%�<<�q�XI���C�z�<�Ҙd�������#Y�)�u�y�<AS�J�=�T� $�I�.y<��F�s�<��AWr� ��?�N���i�<�lX�;�0U)�gN.]��M�<	���l�.LS���u��b@-�J�<G�ӂi�K,o�5W�O5��C�	�)�J� :��\�5�Z`�C�I�Djh4��[�uT���g�RC�UKj��o_,YT @��(|V�B�Ɉ3j�9���B!	��ps��PB�ɨVC�ԉ�H%��p�M��$B�	w�>�Ӡ�Ƙ]hv��ă�7��B�ɑ1���e��#�F���	�+g|�B䉁&_��;3f�0y�.�HQ*�;®B�	�o���9��N������!D'!�DɲUD����)��<��`�!�D�dr|r�� �����*��!�B�uѦb�UxŲ����J�!�$S ���G�L�r��V	�!�䕉�¶��/Li\�q΂K�!�+fw��"��	T��%�N�!��I&!�����!�!�d��R�!��Z'd��ЇQ�jxdW��9�!�D�'�x C�c��[�ف�O�2?�!򤁽�䔃�6'S=8 ��!L!�D�\�khG?�샴��!��٭<dX�ڷi_m\JD��KK;:�!��|����oQ�k��-��I��!��	$U�J4���ùj3j�[�WG�!�� T�Qe�b�8�1��V�Pw"O���B�)�Шp`!ɓ����"O9�"n��7� �Bb�	l��U��"O����ֈ0ʙ*���2�X�0�"O�m˖���Ux�4�_=�[�"O ����*F��YpdN�h&~�r�"O�-�U@"|�)���� �xy�'"Ov� `M�v�`�%s�*	�"O�}���|3"-�@�8��x��"O2�% P�K5+��� `�� ��'�ĝ�E`�;(^�x�'쓀��L�'p����N�byĤGj��R\��0�'�0U{�F62���#�͈E�d�1�'}����U3m%h�p��7�p��ʓe="(iGÄ�nQ��{ �4-Ѕ�3j�R���1Ϊd�dʞ�( ��^���
�ǘ�z���`��#ֺQ�ȓ`;�����Uj��0�b���p���Z�B4��3�"�&U31P\؅����lܣ�Ɓ)p,�	9�H�ȓ^2PD���$/����������o��m��ԵSt�M�@�*��@�ȓ�*y�6�^Q6h0w#� Q��A�8�3,	]�6P�+�+��A��:�Fy1� �7��s�J�2 ��r�4�FFɆq9���@�} �ȓt��M�T"͞
T s�,Y��܄ȓ}SR\2�T��p=��׀D�0��ȓ)����V�,<2�I�Agҹ@��M���L,�G�,�R8���32+����"�K�����k�P&ml����'U����ITHz��)@70ͅȓrp��."iލ���ؠ��ȓap����]� ߒy%� ��5��Z
�&�@q�E����s��ȓrP��g��9,���p70*:.]�ȓ@{\	K��0[����'��2~d�Ɇ�B?�Aۦ�Ǣi��8�B�;xp�ȓ�
�:FN.��=�ы$r���ȓ[w�5"p��"�B	��m�Ux�x��pi�hR��^>��R�]���1�ȓW��rP��*���#6��54�¬�ȓ ����A٢F� �����H�^D�ȓYl�d��*�N��������ʓik����l�Q�|�&�6zQ�C��m�2!#�gR6L ��;�#��^*�B�	1{�,���VI�@��c�|�nB�ɝ
]�$(1�Z�,KL]�c��dB�	�Nw>��yr�kFAߛ}�B�6Hj&�2E�y��9S͛!rC�B��10��*�L�!�����Γu}VB�	(F����%Ü�~�ы���%	�B� �l5Cc�+@�2�#��*!�C䉃 ��tʍ�0�Jd����>b�C�I�>��M;�kR�:���*EoN*@�~C�	�#�b��F��1L%~S�'�*EuzC�I�UB�)�g��h�8c1j��A�>C�IhbE1���&O|-�����*C�I�Oz� W
�<eB�t��ԣ
T�B�I(aJT�;��OW�@�`���^sC䉼crJ0(2b���f/ΉMբB�<WR*�!�NP�� e�ԫH�q6�B䉅h��)D�޼Z6��eE�	�B�%{�MI����Tj��V�-IhB�)� �)�ԩ ���@��#=�bR�"O0tc�F�d�P��"E�0J���R"O����nU?Wwj�� �]�< �C"O̬��D.$��#"�qNH�G"O�H��aٲd�X��Q�Q�^g �Y"O�%�ĦԬb���*`�K�I5VQp#"ON03�o����,�6SI��"O�|B��;?~:�f@'f�@�"O��"X�*�
��`f\/S�a�0"O ��&����@�E\��"O�� �K?����OҰ� �v"O����c<.�p�L�y$�"ON��D�[�N��sьͨN�98�"OB̂$�Z\�5RW�׽,�0�"O�� �32���*�mKt�*��"O�#�M�5>��,A0%.zz!�$�
#�@HG�_�B�6+󂎲!�03������A��Bp��9L!�D�"6o��&!�<q@�����k !�d�3f�ܓ���#>@�I��
�t�!�$����IVjNb��x�d�E� �!��Z)!Q�ؗGp ���M'P!��t�&A���P�ǹV��R !򤉑�b�*� �� Ul�)�#%W!�$ō�~pل�ە7bʬ��j�?uG!�$��z�×�/M`(`w�2t!�Dх�lY�*G�v;(�s0l�+z!�&d��s���-s.����! ��!�$�02�����)�9	v��bq!�dU�@4E˖�ӱ,��E���_!�d\:	1RA*�.�&�*�K�
.W!�U�DC^8ǃݡQʄ��!��*XH!�B�`�(��큿b�RӤ��"N�!�ĈGse�J��m���X�B =l!�dd�4(ǳq�
�d�Rl!�$�:*g��櫐7Az2� ��	�S!�dY�ZϒŠ�ֶtj�P �
O�!�d��X7����b	X5��v�!�ç�ȑ񎒴���K6!�!��?#�D�r�iP/��z� �:3�!��#+6���b��&$�MKՄ�)t!��ɔ|�Ȕ��A`$@��*bu!��)[M<�1N �t%X���"5�!���	���igܕp�A${�!�
�EV��&�_�O�ܩB�f�(k!����*��@$�*0Y��G+.a!�E�u�\��-�z������ )h!�dO~�Fu�!V� |�2�bW�{�!򤞦]9���$�'`V �@�^�p!�dǣ����r&13��)�E �d:!�=����E�`��%	 E^G!�$�$CV*�)H���@ �k!�D�Ig�x��a�%`�e��K� �!��uCR,)`�\9S��8�)�!��2���ա]Eּ#V��9K�!�ݹ\=���P�ցX2~*SA�{�!�d� in�����5�����\�!�^9]�v�� �?0�	#d�[��!�R�<s��ɗ��:R�ȥBf�~�!�Đ�Bb�8�B�=��-A��-u�!��4xJ�����+}�*a�@��5(!�d�f �Gk�� h�g)��Wn!���A�����%F�>� �I!�d�	g��Y��Lr�ji�Ҩĵ<�!�� 2��u�UtU�����&>r���T"O�X!î?N�Ř&�iAt�d"O������aXưS�L��OP`@�"O)C�=�"}1�BK�C�� zE"OHU��W'"�k""��b|��[�"O�ĩ��_/$Yjp8g��bɨ5"OV�闆�*&ډg���?A �:"O�r��R<��e
�2;����"OL�
Ŭ�/<���S�	,9,q�E"Oa�T)f���I�RE J��7"OtQ ���ey<�2�'�4��"O��&Ćb��;2���y��"O�A�猉*,�� �kpع�"O*��'B�ۤ�P�O)ER@! 6"O! @Æ�;s�VJX(%"O�����*D�ݩd�;	���y�"O�$Ц��qJ��j&A Ԥ�i�"OfYHabзc�pHƊ���qL#D���Y::=葎Q�d/��2�3D�l�� jv���E��b�H4.2D�l�R�͖T��Iz
[q&9R4�.D�H�Q�J:U�D�����}$��K�+D� !&`T��<�p�^)Wxh4f7D��R$[% è=�tf�4 �,����3D���5+Ū`��S��Ӌ|���Ee3D�X�A�|������p��t�$D����$(0��Wi�6�����#D��$Y�>E�y`�l�;w�~Q	�j+D�����R9Na�Yxt��*wG\ib6G6D����M��+z�{�.�u�.-s�4D����B�1ؾLm�9���1���c�<�v�X K��9 �1>Cր9�c�<��̔}��ܘaD��<�|�T[�<�eD�6	�$��6��U��X��s�<�V�]W��D	�.y8���c�<!���9&�)��&AI ��5�Jv�<�2�ţ:¤3E!��Bښ�8��t�<a"E�Z!���bKT�~�tC�	0V ���5��b�"U�A�bl�C��?~h �j&�Vl�wM�#7�C�ɛvތ�i2�Q$ � dC ���C��:}�Hr��3n��<2��߮R``C��/+�R�s��1�Fes�o�"=�hB䉓6��]�3L�d���A@Aq4B�	!C��8�Sm���0C��B�	QӜ�兛�slT䳔��R��C�3D�ƨ��#V8u�4���E��C�	t.X�!�o<Q� ����C�5g~��h'ES2�Z�V��B�	�(K>`%4D&-yV�'�B�	�Z,�t;CJ�7H1��[B �/L�B䉐H�����^���a��`��B��;%�@I�O�M�B�)� ���B�Ik"jh{��${Ʊ��@�%�BB�}�l��ծ�.�n��F�QB�ɱrȐj/�,����P��rAA?D�`(uKS�dzډ��IE�`�o9D�p�V��aPR���h�v_x��8D���C�7�^�I�N'P�p$r!g0D��:׍�\���0���h�d�a�"D�����,|
TY�R�	� ]d����?D��1��6�J��%��!�F8�h3D�Ј�N� �����n*�p�,D�lK�/;�l�����!��a9�+D�� ���X�$�K��/@A@���"O���ǘ".a�L;V]�],�!ʃ"O~Ec�lS�4��1�	,��"O����0�� wB�Z� ��"O�D����I.�t�0���|}��"O��:�&�93�r�!���c��l"OT�ꖡKX������J2"O�ĸ��ɱl����Kݍ@B,��"O`ݛ��Ɲ_�`ۀ(�_CPY""O�8�L�?w>���&''  �"O��S��]=3���F����M��"OnA�����P_ )��Fħ>�lR�"O
\���N�ei�Y7��WpZ	�"O���AJfa�e(���Y[�q�A"Op��K=hTB%P`�!I��i�"OXy��G�z`�ٿT�^4��"O�V��J�!f��AM"	�n�<�d$ɰš�&�a0����Ho�<Q�E]4� ����G�u���j�<�P �>2O&( �[�qz<zg�Yc�<�c�
"}*�){w	
7'Ҩ+��`�<���W�nj�� A� h9fQ����g�<�a������@��v�C&��j�<1��	�^y2��K���2Efn�<Q�JB����!	�5� ��w�Si�<����1�J�e� O�
�;0o|�<�1���9e��0��ס��a�x�<9q�޻<8jty��֩R���'��v�<i��űy-l�zNC'd���x��I�<�I|�t �n�TX:��C�<y���t#	�`G�75��8S��G�<1��O�IМ$�'��'�����IB�<qUD�qD�q3�b�9
cvT���H�<��á0�h��U*Y80�\}�2C�G�<Yw��!u�5:�!K�4��˰(�o�<�G,�f��DRSN6-u�1#Q�<�­��t�69����1lGu�<�R,�%}�X�'���@;󏅾�y"k��r.��O�Q��H�qa���y�E�5X����ؔ:����I��y"�R� ���j֘b��y�#�yr�� LE��"V�ԽR,��cI5�y��%'7��`k�w
h��Ua9�yb�͜V��Չ[ ��I�2��y�޲l�8�`����dU!��̽�y�N�4��W(�nwl���C�(�yBJ@�R"���O��`.�c!L��y"��V�`h��A�ZA�@r�)�0�y��]�4��8��ɭR��Z�"/�yG��z�Q'��tt�8R�lC��y�n��E�`2� ����r,���y�AL�_����r�׉�8`(Q�
+�y����
u!�P�D��'�ޕ��^�>���a��C�`���'P��3���k������'��������=��&G�X��d�
�'����H�9�QX,�;��
�'
BQ�Vb�
Hh��	(&�PI
�'5L��s�/|�*�	Ӄ�$#�P�	�'9�y"q�L��~A�ʂm�Ђ	�'���2�] �ư ס��j6����'��A���)Z�� !�̘ь��'�a�Q���P�eѳn�Y�'�� pր��qL�I� I#��r��� ��v�=SnVxI��B�f_n]�T"O8�څ�2r�����cyf��"OR�f�4j6W���(h�U�O�<Y���4s�L�;���DE���YH�<$��G��H�cBйar=�C�<��S� [��A%�U[,��� g�<i���`aV ���  NN��z�<���0\Y�iP!Ȼs���G�x�<Y��1�|z5D�5"��#EGx�<9�'�Yh�ȫЫ��k��ɣa�y�<	�o��y�CA�_����L�q�<��eODhl��3	��B%8u!Bq�<��g]�S��0�	�<&0x{�G�<�u�\�u$�B��J�B�:=��^G�<��O>ܺ������	RƝ��!�A�<o@�k���f�UM�<�S�<Y�ኙ
�-�u�X�|�r�����Z�<�Td�/C��! d��/�d<�p�EW�<	��_�7��X�h <u$f�	U�U�<��L��`��t/F�df���7%�k�<!� ��,ಕ��%��D���A��r�<1�,�K��� bA�a�ębw�l�<��c�d�[���n�\@B0B�r�<��Պfl��	g�]�Y|��
f�<�&�D�0s����F��oJ�u�'�b�<9cH!dչ��ы7Δ�k��E�<�C�G��PHu�H�a��I�<�G
�3x/�q�	7 $��b�B�I�<�" �rE��:͝�/�!"�E�D�<1�h׼j]9D�?�� }�<���
� ���P"j�9���B�<�q�@r���+L�-�܉iF�Y�<)���X	��m�$���1�+ZR�<�PC�&`[���M#h@��Q�<	�l	�b]�D��Ls��RO�<��
C �89�G�:�hE�<�bK&[j�I�۲8����}�<�n+nxޕ���_/4B�l�|�<���Fn�S�)�,�R$�x�<�F2v�u#�X9h�\��fF�m�<1bN� �줒q/�<!@�A`��c�<9�(�
zl{��P9Z��T�I�<���מ`�\��F�A!N��uC�mO�<���!iٴ�p�A(���B���C�<!��"!��I7A� �:Q:���G�<�#"�<UԼꅎÐ�豔dC�<�C1,x�BU�6�thWe�{�<頃 �4XQm�=DR5��z�<� �W���"�ΥKi��!gD�P�<yJ�9=e�� &�Q�6$f��7!D�I@��,1���hR�B�t�j	) �>D�,pAa�t1��TK� �hU��=D�H��"h~�b�$G#-�8u;��=D����U�]�ap��0#�&�'�;D���V�����p���� ٫78D�����W<.g�)S�)\GR���&7D�`Z�	���fM�� ۲�u�	0D���#U]�"%�Q`�0���o.D���F�X(E�$���"�m��ka2D�(y�d�;��m;to[�e��@G%D�DC�ő�]l x��^��R )D���b��eR����˜R[�$
��$D�D!��'�rH��ȇ�&��PrԎ/D�"���NQ��K�d�*��"D�� ��D�ʕ	3Z�� ��k#�� "O|=�c��53��(C�]����#c"Oʁ"'���eS��൩�O����"OZ@�l %������]K�e@`"O�m��B����r���
&h�"O����ȕ�;����o��.���"O��$�j�~�AH[�[��dX�"OhÄ�.�*0Rq!I(Č)ӡ"O�|(A�V.LZPY��	.S�!�"O�D�� $�a8���!�9�"O�Q��N�5^r!4��� �0X@"O�5
ƪ5��8HX�$�N�b"O���ц�(UFI�GS�P����p"O�]���M�\� 4����2���"O搘rA�5%H�&�у���*t"OQ��BQ .!`��� Y�X��CG"OVh+ANp���ʓ1l�%��"Odܸ��&9c�!���ڀRH)p"O�i��� a7���`���M= ��v"O
����;*´�WN]�g74���"O ��L�;C���MA�X.�ش"OĘ���P?Ct0`�,? 6��"O|Q�B��9�<����*G ���"O�%��F�!�vը�D:@���"O����VID"H�j��L���!"Ov9	��[�w�~�w*�+��䊅"Ox���ճ[�j��B*ֵ$|�)C"O�2�EĈ������^f�pJ�"Ohe�Pk

H�f1����=\aN�t"O��-'8Br5��C�v�6�"O(d�wb^3Uj6y�V)����"O��k�(֟)P�"p��h	@W"O�-��EX�xn|�uoݹa�(�"O�X�v%�l�X:2�X�YZ�C"O�pt��/��M�	׏}v���S"O@��sɝ�	�@D�4��we�]�q"O�cD��t8�m�C'֋2^�Q�"ON,��@,ws.�@	�#fV�X��"OD9�@ ٓ/r|!�a�q8R�4"O
��K@
	�V��2��$"�y��"O�t9`鍻vg�A;���>��0"O4Q���4.D���܄L���"O�=ktژC��Р��)9@���"ON ������Bb��"EG0�
�"OġAa�
7$`pM*��E�@�q%"O6�H$��6Y���!HV��1+C"O�D�+f�C��!p}�|ce"O~�ca�؁[�>U��
�Uon$,�yRA��bXi@D\bL�$ʉ�y���$�X�Fd�[�>��2bZ��yb��,�gB�5V&��*"���yBi�����UdXe�%r�'߇�y�� �� ���I�ک� ,Ʈ�y���*}Ϝ�R�ȏT6��&�Q��y"k�D`��j�F��A�`˗�y"U����K��9N,:�	!�y��ڴnxF�j��6�����y���(r�d�2�A7���U��y���&�0<�j�4��]:Վ�'�yҌ;,`T�&H�&}�����ء�y��[�O��a�AR4XH̑�B��y��;p���	��ј[ޚH`Iҝ�yb�
]�VF�[���R d��y�/���\�A�Ou����R�y
� ��"$�NV�����u=M�u"O��ٰ@j��$�EJ�3\Jɩ�"O�x�$���/Pr@�wh�tOV� �"O�P��%/!�DY��C�fC�]�Q"O����.�%:�.	��΍k*�U�T"O �4��.{؍�̖~(���u"ON=���MY��D�6��`�Ш��"On��qk(`�������OEXAxd"Op8J�)|�(����;>�+�"O(5�0���hq�䙄U:��:�"OHA���)���hve[$h`x"O��HE��^�X�j�;q�����"O���n�y$iB�	ʬ�V�p�"O�ųÁ�Y ��
��^�1���!"O�(��ߦ%���sg�$4x��R�"O�)J�kG"	�P��A5Z�h��"O�Y���)��ɛ0��_Rl1�"OV�#���:���%E\BݼD��"O���%-ߓ�h��J;*���$"O2��#㜜fhe�C	�1B��)�"O.��2��z\D�UG�b'�Ȫ�"O`��3L�+O� pL^h7����"O��pd�޵)��U��K*@��0"OF����K#o�ZL�sŇ= Y.���"O�бp�a�b�A��D�.Sh�b"O�АT���`����/{q�P�"OF(IPm��:����BO-sL`��"O�xP�΂�d��f��U�) W"O�be)<��!:�$R�J�!9u"O�����?Ih�@�CZ?S@D�k2"OL�v��!r>�ц`ȁ�~�s�"Od!
�O::�#�/�(Ōi��"O&Q{3.[1���X��U	,�� �"O��$"�|"~i��צ$�r�h!"O H!��V� ����,z�2UC�"O�hׇ֠i���t�[lp�'"O��X��π[\�=�6@l	aahL*�y2�WH6:5��B1|�Q ��ybD3C/u�0��u���#m?�yR�Z�d��E���W�l������yB%D%4;���_/v���Ö�y�V������lH?O1<q(� (�y� �/ ݮ���䚬J� ���<�y��^� 	�D�v/>>l�X�#�J��yB� ]מ��\Es����*	�C䉺Zf�uRR�X%|�х-K!
�C�ɵ4N�PtM2<��XSA��D��B�ɲ7O|�JA�׮��f�k�B�I3*�T E͘M�0!���3N~B��&r�h]�!��zchx���gFB�	 3�� 9��*2��x!�A�W�
B�'D��m��o�uf��(C�.�0C�	�M����Q��Ee�R�K	{C�IhH|�����՘�F�m
�B�ɾAd��O�V�DY�X&�I��'	����Rwv-�$|�j��'k�<xS2;ıc��΅r��i+�'g<���L�4ܝ�!b �3Y#�'��R�T:�(B�N%/qV|R�'�Y*3�	�|V��P�P()����?9X�$��a�p�0H�~/�D��]��	�5 V$z��x���T�N�z���M�ؤbDBB�RX��Z���� D'D��t���0�p��a�RD�#	$D�� ���hT.#�(�H�I�h�Bp"O8	r�KԧN϶����%R����@"O�q�'�mu%��$Q�KG"O�И j��	����Bպ8ڜ��t"O�aP�!D/,�`MI���.���"O18�-N�x����D�O���"OB�I7���tД�0v+�3:Px'"Od|�Du�2��������"O\�5�]R�2l�@�_�ʨё"O��t���wp�޹N�>�� "O*Ecy#h�S�
\}�Е��"O���g�7�
�[@��m�.�0�"O��
�@����@AA�q��m�r"O��B���b���aϪ��$Ѳ"O��*��Q"7)H�C�ԝyp�y�"O(�����&wtؖ*|I2F"O�tR�+SYU�����!���4"O��iv�PT�>�I"g�#��)�"OT����Ne���r� P��Mh"O~tAf�'&�������>���S"OJ��a��)�Pڴ�I�pvY4"O����d�x���T� 7L�4"O���2CJ�K�6��(�+&��ʐ"O�z���$#���WɅ	#j��3"OZQ�t"�&O@|���]:Ωxp"O�)��y�@z�J��Vﶭ��"O�$�@��?EٺB#������W"OĐb�#�#y���s��'tR�"ORUsR[�#�v嘖�A�&���z�"O�h� ��u���R�Bi��:�"O���A���?��ŒK]� `"O0���(&����'���L܍s�"O�8 
�Y��l�,2`
(E"Of��P萴AF�ܳ����]�Ę�"Ol�R�ޒT�@�h�6����T"O �y&�?��b�س`m\�j"O���4��0!��H��ڵ_�,��"O���b�Q��q�w�:'dz���"OrQ3��$���kؓS=�\��"O4$jPFY�JQ5;���X���%"O᩷��B׸dAa�X�s8���u"OA�W@�t �|#%o636�:�"O���$j���x]�Tn�+'x�Z�"O@L�eJ4pTXҡ�&}�4��v"OV���5#-��cԗ..�-�"Oʽ��/�d�l����D�eXLj�"ONEs3��ePl�jg�۪�����"O�x��Q�S�a;�C��P�ⱃ"O.���V�:��d`\L&����"O4HXsl�+!U>q�r���5�.7"O�8���O"N��EJ�->T]�R"O�̻!��W�b�Ƞ��?#�!j�"O��	����4�@�	�%��"O,i��F"�|���O�x�#�"Ob	XF��9R���`H�S�"O|��� ݧ
7�����ٓO=���"O�Y)�ύ�-�(kGd���<�C"O��H���<$j�ī�עf�3�"O.��p�C%\�RDB����XV"�{�"O��a�����Br�Ğ3�.�+"O%�#�+s�0���R�Hmٔ"O�A�FӪc�ƭا.H�!��e�5"O��woA�n���#I��N��1"O �I��ׇ}[� S%�ԚOu���"O� <���QLW�|8��+a��|@f"O�Bt���k:��JJgʠ"O�q0��.� ȩ�H�.s�r��$"O��e�	 D5ܤZ���5:��G"O�I�&gP`�$�7.Y%Kz <��"OrMa����s�Z<E&˪Xju��"O����h���$�^�=gΩ	�"O�@���@�,iI�G�לi)���"Or�{ +�4Q����R��ѹF"Oj�+p&�5xPީx.,`�B=(�"O��j�M�h4 ��
A�Jz�1"O�!	ff�
&���ٱ��t�Ф��"O4�;��׆���B3����p"OΉk1m^[�}��O/�$�F"OִQ��W���q��ʝqu��2"O.q)P/ ^J��w�ʧ3YB�#�"O�I�V%�<G�Њ�-@
�F݂�"Of8#�IO�fLse�J�Vq�� �"O�͢��ǙIŊ��g���2}�$""O�ɛs��L��Eys�H�pg����"O|[%LϫH�d=S�Ƈ7�|�&"O���A��J��D������ �"O��6�J�y��p�gÎԠ4g"O��j K�3�j����;m��;7"O`��`���$�R}8�+U�T��0"O"m1�l@5k2�Yh���V �"O~��f������æ�ȴ��"O����ҙX��  �v�D"O� �q��Be0i�oT\�ݸD"OfpA#�|�J=R��A�YV !Y"O�j���>)���(�.+U�Z�"O��J"6Z�|����Ie����"O��D��ug�%z�M�>�Vy��"O5ȁ�+a� xs._��jIۢ"Ob�8�R�ВA�핡(},t[�"O<(�K!����TM�1N	*�"OJm �`�"i��ܫ�I�#�f��"O41:֊��'oD����?�z���"Oh��"��C�R��N�q�"Ox-�!Fb�m���Pf��t@\�<q�!�\o)���-��
dGM}�<��"���R� Í-F�*".`�<�	�?��jD�b�rl��w�<��P��l�pJF"@�jɡ��QH�<)�Jď�HE�я	�sr��P��[�<��m��q.�0/	�1 !XS�<94�ėn>4<k��V'�1�B�v�<a4� �nϼ�yШN	j�.��N�w�<�g�ئXDҰ"󇏐)�|�5a[�<q`\�@�D�*�c�5'3���!�U�<�!,|n���
��on��c��Q�<q$�v���ڃd�
�������X�<����-�u�BH�t]�El�<a�c�"݋#��T��jS
�l�<�֦�Z�`�����W�D ��DPi�<����i�b�s�A�N�X�#4"�g�<���s��טB���{#�g�<�� �6B'����V�D����^�<�
LHvhx�V$B3�<���S�<�pi�p ��s��A�7?N�S0��T�<G䌈?��j���C똭���S�<AR��uV0;g,��ZHJF�<qB��r�X����`z�`4bJ�<I�kOl��A6(��c*D@�	\�<� �#6ꆧs@�h��KK�68�a�"Of�ʰ����A� W���X��"O����%	;�y�@�ې�d1�"O"�V�� ��M)C���S�j��"O"�JW�����4ף4�d`e"O���5�O01b.T��cQ!	�\�W"O�h��*%���ӡW�=Ϟ}k "Op����^(s��˃n�Gi
�R"O��vK�?}�p��L�0cF	�F"O�0��ك/��Mj����Kc� a�"O^�h����=l4Wa/4Ot��2"O�P���g�Ȫ��֠79ft�"Oz-��J��G�r5-�>	|��"O���B��8۴e[�̞Q��1`v"O��B��LȌA�	��T��y��"O��z�c�E-<l)t��B�$�"O�͛=_a�9�rk�Hr$��"O�u��H
<V*�[!*ɜ1Vs7"OF�ŊTx�������-�ڄy�'��$���A85��{2�H�x�pz�'odE��gGT�r�H���m!X��'�h�{�
�;D�	�1AJ/i ��'ID��s�@-V���`�<6϶�X�'pް b ��vڒ\�g�_�
��'���b��2$u���엟M���
�'�bX�._;6DгvbޘO�<��
�'������)B|+G� @�BLy
�'�� !��
,�F�Z*�
�2
�'q��:���\e��	�"�$p`
�' �5�7�:/-��eݫc|�ո	�'�V�×-�$����;���KK�<�Ui�?5@�!��8�|�2'�H�<ɲ���D�����R�B�C�E�<A@��2.���B�yI����i�\�<��E_Ba1E�/SST��V�<Q�� ���XǯBT?l�zE�WO�<��T�&ք|��
�m� T���J�<��8I!ܵ�a��/K5
��Z]�<��@)g��q���V?Dd��S`Y�<YEb��i�P��geޑJq4����EW�<Y�b�$_L �Юǲ.�� #��}�<9d�D51�,q@m
.o 9D��x�<y��ޣS�FE;��|z�q�GI�<Q�C�.Р���Q�q�E+�E�<ѳ�_:h�����"7h8*�%�w�<�1g̝~qh��f^� ���9W� p�<�gO9V���b���*������w�<�֯م7�B�s1�õr��M!գ�z�<1�M��<%�AbX5zN
A	��v�<�7��;^��c���5P���r�<�c�\/g�@𷁃�J�NQ0��r�<�����CIP�@)=�4�Cm�<I�+$�\q�����E�6�K�-�R�<�TQʜY�̟.7U-)CAj�<�!�
d�,�څlϓnX�� ��Ai�<Y獃[�m0p/˫}/p�Q�_g�<����:`E܌���+T� Ҏ^g�<��g�5;��aF��jC��\�<�fLC�������aܸ��@Q�<d]=�|�c��w�1SeGM�<�&eЉI9�|r2�M<7;���!JT@�<��D�c��U�^��ԦGy�<����qxV�2rJ�c��I�<ip��u���x�R9���7��A�<� F��F���+�lP0��;	�h��"O��j�n�
��# h��s���@A"O�@�$�yI���bGGe�L��"ON�`���0@�[�ݹL���"O���TE�T0pf_e2h��"O��v�5Ovp��E�!W {�"OZو.ںm���:�Jŀh�j�R�"O��IG���`z��aD	��E��h�A"OB�@ׁJ�m�4�K ��
�Li�"O�k`n�S,TiS���4*_P��#"O�	B�D�dF��CO
����"�"O9P�dКw��Iюݱ�"O�H�WHŸ�DJ�+Ѝ"P
���"O~p��cݴ f��34���δ�"O��A���
Fe�d3�\�Bh�iC�"O^!����"L�S��.=n�sW"O�%�䈖�-� ����@�6"OD��%ĝs֨��Զ��8"Oer@�2w���G �Ҷ0 �"O�Ꮡ�H.A��i[�h���ۥ"O����l^'P��˗�� eo�l�"O�0���`����oW\P`A�"ON��l!\�L1��L	:�y(6"Om(���b?�!V�Ѝ,$y�"OP�Rr���5g �"�DZ�R�2b"Oj��!��
Y�+T�ٗ2��k4"O����X�{d�+#�׍]���;u"O\���σ$I ��i֊�1�~܊�"O J��G�Sh�!����&�t�I�"O(A��$8�!�0�G$�(ݚB"Oh����CDy8��0k��R�"O84�D��$��ҡ�6��X��"O���k7^�2xJǠJ�iu����"Or�R���4#��\sq�~�5Ns!�d-��%�0	��{��|�dB?!� �	ǃ.[�\��R�X;%�!�d�-p���*�	C��@2��?c!���>iij��$l� Ka!��7(�j��vfĿS�ν�4 $?!��n첉�拟�nh9�h��!�D�m6X�U�BV�V]���غ�!�uƾ��+�sb� ����!�
�mh�թ�e� Q��A�f͖Y�!�$
��ȋ'͂$��T�&@�,0�!�D�#E�Y�$���\��e�#�͕P�!���r��ߤ6l��	u�Ϙe�!�^2-��@�!+�IW�	S�O��q !�d�Q�d|���?��5�^�!C!��ߝ�>�*Ӭ���2ДmҘ>,!򄌑5+V@��D�U;<8Ы\��!���*��qb�,99�����T"O!��V��}c ͝M!&��iMm9!��u��E;v�2`�{��Ơs
!�dK>\���C �N�g���CJ� �!�94V���%RL���B�D!��)$�B����!bA�t#���0e%!��P!%����&�&FE� r�&�!�D_4�l�j8��M`F�Ҧ�!�dH�W"�(���W9�Z3��N�"�!�$�!D, 2lKqP@X��\T�!��̽i�i�B,Im�@�,F
um!�����NF�,iJ��B,J4�!�d�
4��1�����Z	�R�Z�j!����̝�qF�<[S�	�BON�\�!�� ��N��M�;â��Tu�'"O~���'�8	����BY,��"O�mA JK��&�#����V�f�Q�"O�	vOE�Xe��1;ך�)�"OJ�
�`P����	�3�:)��"O�ٓ���PAj�ruI}�\4��"O��k��\�1�������%�t"Ob�U�S~���W �h�����"O��PfbK/8�x�%��9����"O�S��8���ć+���p"O�cl2'�Ո�ܪ^�`��"OZ����Z`�ҤK�{~r�
F"OT�#��D5ot\أ��5N��p�"O.�@$��1�pݰp&�6C%�r�"Oj)�jJ-��iJ��жb
��R"O^1P�Q�	!,c�&�I ��9#"OĨB��S�tL�$��-�Ҥ)�"Otu��ژ�BP ���0b���xA"O���@&�f�*Ah"+Ґ{�V`��"O�)R�A�NK�]Z�i/U�8�"O2�cw�P�gb�rfi	"T:��u"O:��� 
:�`�Ҡ%S?WM���"OVEz�a^s�����)�"UK�"Oꬃra0iq����M�T��D'"Ov�K��� �r��2��$:�!�W"O���KQ,=��i��]�(9FXJ�"O5a��F�f�>�����;G.�l@3"O4�E�?(N� 
��v��8�"OF�C�!B�K���k��H3�$��"O��L�<�����	$(=F�ط"Oj8�JO4x��F�۶z&0�Ȁ"OmI����Z�^=�RMF�"O��N�2�(�g�ڇ�P�P"O
h�1���b��ۖu�B�c�"OZ4�F�	b�"�*Z(9w4�b"O�u�1�
.��Ui�iW�uJ�:&"O��g���ހ0�ciQ&f�u�5"O�b�To��#��K'��8H�"O��A��8ʄ!*Ë3ꖝ�"Of�F�$��l)D��O��x "O �[U�F�Z���$]�Tz��""O���m�C�D�� �4uŜ4�"Ov�(��8��0���^�:d�'"Oऐe�-��URu&ґx5�2p"O�m����>Aaf�2P���q"O�.ќ[�F���"z��3�"O�"v�eW�����>5"��"O��zǅ$1Fh��A�y�N��v"OL�^�3�8�1d�F�\����"O���L�dxST�>h��i�"O��	A��+��%��
ܾq����w"O���$��)�jk�'[��<Ba"Od�E��=x�|�&H�/i�J�c"Oִ���TYqF\�F��X�"O�Q��Z^~���Y�V�l)Q"O�$
���,|0���E�UP�"Or@01����S���Xi��r�"O�H�e��R�HųcD�kkd��"Of����@�Ru�X*��ҩ}a0�"O@�q�
��_����h���`�"O&����3i	�A)�!����C"OTe�5	�6�<��&ҫ=�
嫕"O�4��K�.��&��q��5��"O����P���L�E� ��=�#"O� NE�&�΁7R0�q��?�b�hF"O�@�e�:��!���g�~�"Oj�w��+9��%���	�Х��"O0����	�%�"(8�NE�]ͦ�:�"O<ܺ�̅�8��]	R.Y0��*&"O�$�eO�Z&y��.��YW�q��"O���Z�~t������[��bq"O�[�*&$�~��A�A2ap"Oh� ��?h{D`�nY��ؐ��"OX�.':��`�.6�lD�E"O\��AK(�$*�fɧ<��R�"Otɣ�e�[p<����ͺ��"Otw���!Ȗ�Kq�(v� ���"O:���\�825 vLy�Z��"OV�2$-P�A����]+l@�cW"O ��fj�0���VH�n��`�"Oƌ����Sm�9��Y�y�Q#�"O��
ޠL��(�J/+gxi��"O�)*"(
�B�$���f՞���q"ORyxG��,P�8�)�˖�>;""O����`��s���ӫΤȀ��"O���'^0l $�R됿oJ�r"OȨh�	�0tHI)p��(4!l��"O�	�I��R�� ��y���"O��g���C{�X:qJ�x�$T�@"O,� �U�ndsvh0`���B"O��+VC� ���� �@��,�s�"O\$�E��R�<�G�=L�u��"OԃbM�	�D��&^2�$Q"OT,�A��E�t�dW�r
jii�"O�mY��۩dn�ʆ%�	T�\Y�"O� �	�e���Iwf4��P�r"OH-8�AV<V�@3�ͽ,�z* "O갈�����̫R
��/߄�q�"O��c�K�j ��W�
�p}��"O\�bLC&\����U`s�q�w"O�)�Rߺ�{��Qe�\��"O2]��$Q�f���̮����"O��U�>�  ����B���"O�1,�oΡ�"EN8B��
d"O��$�U�]�1r��gZ�7"O.}�qHT;zG<l �T�=`�H�F"OB����c2 %��$ѴzN��"O����I^�*ԠI�&��Aت��q"O��ె��G�H�`��F'^����"O6ĂF��6�в�l[���8
&"O|yZ`ꏱ=��Q�k�,�\�`�"OT!��oܦ>�H���\�8��d"O��B�i&zq�E P�jĠd"OVl��
Ͽ(h�Y7בW�Q6"O�yR�M
��Ї�D�bgl��"O�PC���+(�Z��E!fd��v"OT�ڕiC� ��y+� ��z&|x"O �I�Ĕ�<��K`S	
y��"O`�2�瞽PUԭO���*�Ѧ"O\)���ڮ;o�	�%D��0�e"Ox�J�.�yKFc7|�x% �"O��t㙀xw>AZ��[\I���"OFHH�� :>*)�����HB쵑G"O�9"�G�������%!6bEB�"O�0��@X!,y�ۇF۟kSF���"O.O(t "D���#8(l�p"Oڽ(SH����y�zXE�"Ob8��Es}��c��^�v����&"O� �-���\�#rp9��xh
��6"O�4����)~n`��p�:q��UT"O6,p��<m`a3/�D�P⦀��6��#�'0FH(�a�fecw����(9
�'U2@�u�1H�N�*�n^	Y5�8	�'�0���˒�V�,R��%�X���'���r��F�{�$�6 ��c!Ɣ:�'�|�Rd��u&�ʰe� �'����c	�}�*�[�*�Yu~X��'������@� 4�m �O{�|�'j�;f�K�q�2%Ac/�*�N��'�<)Q$�SS��,(�"�	�f$�'!��B�<	��c#Ǌ����	�'J�����6�$P	� �^���'�>�J�(ûm��H�E���d��
�'��M���XWBp	a�	�Zo�
�'��P�	��L� ��^b��j�'ؖ�y&�':���С�J=�')d���Dխ[��%��V�|A��'�Tp��풉[0bl��E�~�c�'Զ�3IC��*����:h#�a;�'���ޛ?��4��e��g��c�'�����M��qr���Mڿg�U��'�f�a�j-J?~��'���M�z��'٪� Θ�:��	1�K��;��$k�'݆���hÛw��X!4b;�D@M>)$"�;�@�<�}Z�`�5DJ�Z�-H6g����ǌ�e�<��&�";����QCM
?���PM�:kT%&�T�!��������)�g��!�a���8�H���y���Br�O�	x�+&�Úx��"��/'������x����JּY�Z��oAy��1��.O���
��|��;��h}�(˒r�(��M-%�A��'���y���:1�8��	${<�Fm]���$T&"v�̹��Z�qښ���S�� �`E�N��<dJb��"�@B��.6���r	V�}�@�oIi�F�2�ϯ(���̴S��l�%����-Lw��:�O,kWRpq�T�:�}b�Խ8����GJ(��3����	��Q���.G\��P��W�y��x>��J5*�K8�Lz2ORy�uEz���<ot�*��@�P8	��j��>��	O�o������-�l�#��RF!��.0�����]<�����{ܘ��@C�?j4��ա*86���M�/�H�׍�R�4�k����t��G8�y��2xz�0�2����|A5f�D����狂/��C���Ph�L0�Ox� Dy���F�����HF��7�ٖ��=���8x�I�Њ
pd��)A#C��1!#�`P�Z���~�
D��s8��P/�&O��@����<H>�LX��;����]b��H�J��r)B��n���N�?}��iI9:d�����![؀��+6D��9�!L]n��@M���MI�E��?�8��bk̂���JbTVL�3,#�'�y'/K3`^�E
�eчa�B]��C��y�g�,l��|ar��ؼq. h�U]�Xd1�pa�u+f(�����𡰆�a"�j� �
<�zr�G��
X�dÌ ^�Z4JE,�!�c��-br����B�JH����>�<��d�Nyniy�/�a@�(y� �"�qO��I�G����H���
z��4{�$��~i��L�e�c��]��`�0�R�S9�H���Pߖ��/�+Q�aK4��q�>Hj%����܁j���5B:����"�Sj�����LuY�`�T=j�R�m��3�!�Vj}4!V�Ւ.�ɠ���rxq��gS�e�B�@ݏl��eCg�h{:I��H�y�,��#�
dg�ap��Q�z��Y�yʈ�u�$z���cN9E��5�Gj�9X��+#ǄO3��꛲{�����9(P�6���]���TkZ5�qO�]�E�N�^rr����5t��f��Y�����[\��oD:��ڴ���A�ȓ#�l�E"
b:l���o�D8�� 2�G"Z/�x×[��Mq�"��rx��w��<��%����Qc�\�$Kx�	�'	���3�]#4�\�C2���+�ʨ9��<�9��P�D'��W�[hc؄K�G��hOr!�̑�Z�8��xQ�ɛ��'`|�p�
�z���z��9� �UZ�J��gCة2��_)?7f�K�LZ���a�'���QC�(a����լ�+dZ.ݩ��,�$9���C���S�,U�������^�d����\�j��ԦW&$ C�	�aD��∕8cpBQKaR84�V��,�P�+6g4?E��'z�)�K�F��t��U ��
�'�����^�	;Ԅ�4Q0���'�ʘ�RX�'����͋^�|��*S�m����)[�q�!��85��Sa���B��ţ'.��7�!�d�����g��5lت)[coD/Vh!�D���`hX���	��h�ᓾ5\!�dT!<�F(3�@ 8��	{��רlI!�xs�谕KO�,�P��f��V�`B��7����D�@a[��(TB䉽H4�P']+P�0�i ˜)XB��-P�4�Cj
�T �f�QP0B�I�M<l�*�ŗ�,��׷rB䉖\��}+�m��AFI��.ɷi4B�	2m�����ПK&`rq
/.�^B�ɿg�|��+.a~��R�IW�'��C�	�9��1೯T=m����W71^�C��|܀4��Մ4ʹ�XbgX&�hC��$/��!���4p��]�&
YqnC��n��j��:q�b	��GR<D�4C�ɍ�\B�D�0,����KE�t�,C��"5�-��E�(&�@��;l�C�I�*��aG�P�E���Yr��!M�B��3A��Q�H�!)������Ɍ<��B�I�|��BVoޥ�M �Α�k�]�ȓ
Y��AE�K�"��',���FQ�+�k�b�b��@ߨz~�ȓ$���R ˈ_ِ��vɤ%�e�ȓ_�\Wa�9�z���G�-8�\��0�V�R�GU�e}�XBv�(Il��	z��tH��T�9*g��^����ȓ<o-�q)��x�Q��#	�`
؆���zv��M���RB���D:r�cN>Y
�b��%�`@;�z�е�HuɆ�	�<��,D���`�>��Y�0@Qo�<�w ԍ.6~�q2�@w������W�'5?%�7�-e����c�;I\��U�'D�<�`V%]��xdꓣ��tz5d�<���eц5:ĥ�5@%�p�Ňċi�B䉭9;(�y����� �C��$��O�����q���f^RU�e`��vY!���.�r'�G��C��<\!�أH
��`�K�-%�Q�b7#!��}��4���E�c vy+�c!�d�hm �'Tl_�(�$��D!��:I0l�ȇ�;ݎ5�(�-�!��ʰ=�L�s���'����E%^�!�V#,F,���X�3�VY���^�!�$D."�iG�1���8�N8Yz!�$�.Uq@���R7�~(���T!���k���Ӓʕ�4���
�@YQ!��yA~ԙ����0�D)FE!�\"*������]�KdpH��R!�O����E�B�7����.#J!�dƿ/겑WmI�%���a2 !�$
eX@5�0ѹ[��%Kt�@ I$!��60IAI-h��	�DL�<'!��q����g�=E�Rqu�0�!�d=[�P9@�R*i�Q$J�6yW!�d�K��YI�G��EF4D���4d!�$�
`>�M:4�7!$�IAƎ@!�� h,��n�� ��i����4��X�"OayҢ�02�� W㐙W�|=3�"O �sff�`�h�8�(��Lpu/��gg�%�=����Ob���5-	dh$쇨S$\�H�"Ob�떉�xҸ}� a�%(^(��-��o��d��[�a|�Ѱn�L%��ݏ�h�b����<����x��Z�]x7� 6w� �a,"8Lp(y���V�!�$�c��;�+�0V̨z�D?3ˉ'a��I� ə|c�q �Q�q&Q>y�	���U�A)� Lb�l�5i(D����74��Ba���U?z0b�e� i+>`s��ެ��"d\zb?OxlANӥ~����.v��:A
O4�8�HV��Rh�q�<�^�[�i�%�n�Aq*��O^ы��9�0=�b�K/���I�`E&LH���SI8�|�ׇ�"	�֏N�O#�����'��1�/͍��@�Џ	�*!��+C����T:0��"ՎۺO��I�uc=�]���TH�)G���貫4�S�P ۧE��*I��-c��B�I�v����ՙ!���1&��&L�8����l�N�1���b��i)R�)��_��/h
diŇ�]��T)2cY*BB���in���T�2KI�>���	]�<�y �D�/���ë�qx��[	@?��q������x��0OX��� ��I���Gl�8��9�4`���JE	`������!
��!��B�ɜC�.�J�f�)L�傠ՠ.I��S�>9�ڨGP����ߧ[��`9����$K �����?o|��ԩ֦�y�aPzN�T�&��b;�YLX���"i8�[��mA���Q^p�|�I>b@X+e����	�2 Qa0GZE<B Ho��1Nզw#�����Q�j಄�Yv�BA*�b�-,���y�|}R�*C"Y�,ѕ���~>r܄�	+�nQ83d� *`����޺^�,�!��[�@�>́VB�'8E���"O�E� ��q����!a�48
}Hd�>)�#¯'n~4��E0kP
�	5�'�`ň'���h�=1�������h�L=y@팋g��SA������)��Ĩ�Af�O�-H���^�g�	�V��7��0Y���w�R ӰB�2�
ś.$͔Q��Ե	H��#�,T��j���:lNY���`� ��p�݈Xt�H�1��g��ĝ�Yw�X�qߍdy	޴n�|\8�&��,AI���4������ �$
/E�`���F�� ��=aRc�}�X5 !�YD���
'u���늆J�����V�,�+"��8��QxU�Ƹ��%j��R<"#qO�}�#q�E�QP�}�,�'�F��ͅ�x����$�.L(t"��F��\�ȓ���@6M�Z�.���/:�����3&Xr �ׄ3��l#��P����E��Y$ԖxH�r� `�^1�ȓW4��feE�:r���q�$��ȓg`�L�D���'|�8��ō1H�\�ȓd!��u(+'I�Y��I�J@%�ȓ|���('@��P�bir��Ŏ(�zm�ȓu�ԋ���3
%��G��|x@h�ȓ �(8Cq�K�"��@H�cJ"dS\��ȓm�@]"%�Z" ���A� O�PFd�ȓ	�*��� O�F ��+U`��؄ȓ��ّ'%�='Z&(�ge
2g� �ȓG8�`���jh�����9k��D��3\z	1T	]=V�t)���"�r0��o�a�f�1
״�x�I�5�I��E�AC��T"x�~��v�K�Fä���Iy<ա7j�~�+�,�Z�"O�Uq���k&pЃ�9P���"O�,;��XjE��O��P��"O��dĊ?�Xy� c��R�"O��y�$#d��́r
*	��2A"O����#��ib��#M�V� B"O�0��l�")a����ԦG�ܰ��"O�h��JX��DP�Ɗo�t��w"O� ��3N�� (B��.��	�3"Ob��!�F���3�$V	q��}��"O��:�HS>Ov���B��6��@{A"O�f�èq*U��"Iab6"O��B��D�e����i,P�I�"O~IqQ)�h�����
r��"O��F��k�!�W�AV#�S�"O��0'�8۞ �U�\c"O��Ɍ�$*"�Ҕ�(t��8e"ObQ�ƀ�0Al,��U��Nm0"O\�9�
�?I�X=p$�<%�,�a�"O�!�BK�< �y����t��w"O�i+�N8v��a��(�+JF���"O�<���>?�$I���ų�8�"O&�+� ��z��J��;F�fȸ!"O�2��E�����IѦ(� P�"O�C+H�]�(�;ʂ,�"OR�p�-y�d񐗍H;x^|Q��"O��14��r�
�sBlL9.2���"O>$J��*Kx&���+B,'�l�U"O��y��l{��4
Cw���6"O�9�#�֛w�M�6-� Fm.C�"Ol�9P��8.� SL	�T�,r"O:e�#n�1y�✋��]�*���"OxA�a�C���
�%��^h�r"O�gF_���w���u"!Pu"O�L��&�7����Q�E:qT��"O�UЁ!�T֮�`��? mJ49�"O��a�/C�7�L�
�� z�J�p"OB�:!��(W�"���Nݣo�iY�|�n]�n�mQ�y���aȚRm@e��Dެ<��0L���y��0�-0��\
0�p�n��4���K<�BO�%m���'����׹ay�9��M
�s�8�	�'��\�e�%��!8Dhϗ4�8P�lS�Y rI`�߂��>�' d�HQ�r�ָ#eFy(��CO�(�JB ��SJ����J)�X�b�w�p�rC��	=�!��ɸC���Z����p���2���s?\B�� �4�8Z�0�M�M�d ��\���rV5.C��>��0;g-H&
r�����t$���!O2r����9����b+��$Ԉ2)D�8 	�.2A�h��N�}�+��LJ��8?.nA��j	$J!�x�� @Ȇ��3b���P��7�<�nIS�ܰfdJ�uI�EFz�MR�pp2ǄI+PaF<k�EK�&���"��\�3v����%�!���8� ��4k�� ��Q�Ƶ�p��S���L�
03� ��0zps�χ��H�'J�:MtȺ�ֱ/�<l�����y""�*p�<�q�f[�!��k�*�e/D�:g(�m�y"b@�>r���!�O�:�EyR̀�^:�����ݜ$���ȥ�@��=A���_� ����Zv��@���e:y�#� P=���	��P0&G8����`�&��2�J�cڞ��T�(���|��8q�# �&+Z�õ@T�=ͦ�>Og���+C�tp�-��RͲu�wl!� �B0t$��#G/0T$`q�E�q�<4+�b	�t��5;��Ôs[p2���kޡ���X ?{�9b䞟7Y�t�&D�LP,�y堈:�\�>s����ǈ�@�ڡ�.K*u���獊=t�֝0un�Gy��͆C�n�S�H�nD�%���>�p=!�*��f�dmV/S�1���#Z4DH1𡕁s@8tb�*��i2�qD�|J��XG���eN*1=z0������'<�YU���B"O��(|L��a��\4��o84d)��ڇZ�122a��Ud$C�ɍ|���!��<n�d	�ʝX1���i��d~��KƉ'����O�~���d�țw���j��ؓR�t���[�l��
�'������I����v���c�P[�)^~
���Lh�Q�!L6s����w!@K�'*�$�RLU���SfHHYZ>Q�ד2ŘZ"�WH[���"��t�-���B�T�ta��%N�t���w\�" S�'�^��ċ��n��0Z.�6�p�؍{�I��x1Xܢ&$X'.P۷�� t�"���ä?Q�Z�Dɻ���?@b��W�4D�� <�yA+Z�6��lB������E(C����3��J$@x�}� kI\�:��2�+pޅ�	D>wh P��eIwni��0D�p��ey<j�!�|�[-�6z_q���#2lp W��q���W�'���a��[�� �W��_�����e�b����Z}�i��M-1���7�/�pd�d�.1k��bP㞌~aa~"nR7}<a%T�59��!�	�	��'�>��\�!h�l�Fʨ'iv4�K?����=*�!a�
X�.]���ybA
�X/jm�iԛ%�ԍ󤃙�$�\��"և3�@�I�O?�IS����/�/�>�	Ƃ�p��B�	2��c�(Z7>t���v�j�I�p�D٪��K��p=��+�.i�x{ DO�#+�]�f��w�<���K���7��0A_� ��&�q�<Qe"��Ri2�y`�C�b^��c-CZ�<Q��P:7H1 #�Χ@�^U�C�Z�<IP�S
|�P80�T432��s�bEP�<IS��7*t� DD@�1��pK�QN�<����&��E����1Y�&i!MON�<���5y���2@\F����Cc�O�<�q��}��g%K�_Ex�F�c�<��ŗ9d�ȅ0�nҸ,$�E�X�<�#�	5�(�	�C�x���L�T�<Y�ˈ�eDP��4R��I�dD�<iV Qq��i��
݈XY��3([�<I 	<#�5:�j�2&,"���@�j�<�7h���x��Z*X˜�)u��e�<���T��l�S��*{�<צ�_�<9B�P�}T4�Z>l�FI�@��c�<�o��%���ЬE�H}��f`�<YG�T�LeV٠���}���g(h�<ٱ�5=�HQW�I�So���S�f�<�Q��U�Y�)P)���F��{�<�#I\v�@�� ğ�6Y��)3GN}�<�/U�:��Y�4�ڹC^ �$z�<����SS����H-ᕉ�c�<��Ju�lm�T� PT���E_�<a�Hӟ@��A�ǁa��83�_Z�<�@͑�ZnI����9��`@P�y�<I�FQ�M�0�K�"��4���	{�<B
T2��3v�M	U-v��� �{�<���@Bq�VH�:.�k7�q�<)a�������#��6�n�{5�WF�<�!\�3�|Pj��0�:�ك�I@�<Y�c�6�� J��_H��Ѷ#�<ybHd�zD���A����+��O]�<���J���v�@1=�R�	�fLZ�<��
6c҆m�OZ�J��0�
T�<q )�!^.�҄̓*k���AV�<�P�O�Q[���#%فl�8�:t�Q�<	BVcp�PU�O�p*j�Z�!�R�<��.I=)��g�?0�NeR��YN�<)��+����@a@�J����v#�c�<�u��>�4���ʁ�`-ji8��NP�<���1!&�k��E3o��ԥ�F�<�3��y�6�q2��5L��)UNG�<a"LֹQr(@��O\��y�MRG�<E�b��@�G�W� �pծk�<�G�	�N<�%BS��yG
�\�<��n�u���� �֌ PѫHf�<�'��uOLE4�C�bRtZ�#�b�<�S�G��6 )�jx}hPX6��A�<)��V�m���Q�
fr�ID#�B�<��D
�(��E[�DK�,�dx���A|�<!6�2n]Y�i�2 ��r�{�<��.ҷ�*��`A.Bդݰ����<� Leꐠ_�`��C��S�����"O�d��_
c)� ��H͌[����"O�dYF�¹.�<�� @�]����A"O�ID �2慲q/�%iw�Ő0"O��kC�p7#C�P�q� )!�Ȓ��6K_5E|��c��H	!�䀲W�´+��O1,�4,�e�!�D��mFT�r�$M܆M@�N[� �!�۴?�i�7�7/@����.!�>l&�X�3@�pg�ݣh!��M9Qf��A�L>��Ԃ4
Ĝ;�!�D�zj��#�nZQ�eɥ鐁;7!��S$LЅK���	��XY&'��f*!�D̙g���Q��
e�X����T�J*!�D^	3�u�R ҙe�f��M<g!���H�NԘ��z�g�&�!�.;�	p��S�D,�I��!��<`��Y2Ʃ�x���:�5	!�d�|�|�!��	)4	��S +�!�F�B�l��cӾ]�P�yS�Ŵo�!�=EĀ�����Xr,\;�lC-D!���:~̠u��-tb�푲aA�!���6�T0�IETv����.�!򤛮fe �4ϛmBE{�5�!�dN�$� ��7�`6�Z�A?>�!�D�ܙ��Ǒq���g�=�!��ɤ$�0����,R,�AB��(=�!�DD1B���� L�4�3kT z!�$������.˧>�3#���1!�Ě�n'�����L3?.Q�1Ɖ4&�!�d�4�%ʳv Kå�y!�E� g�D! �,t(`�J^&i!�䉨I5�``�*çv�"�:�
T�lV!��U��4ѐ-\aX�JgI�(jN!�X�'�e��iܓ?t��.�v-!��L&�t���P:�d�ʑ�عi	!�d�(=f��+�6,����g�D�q�!�$��pb��B̾CZ�`�����3�!�䂖W ��q�H�'�:����'�!�$Ć�x%����b��tsGR58�!�~ lh��Պ[1nih��{!��!Rh�V�֩�&Z'�E�({!���
b0t	���cI��;^�8$S
�'	@���H$4
裠�B�`���Y
�'�������2,�iA�Em��S	�'�yYoW�=ݼ�!��ɞ5P���'-�T2E���1��� O�6D~���'�Ģ.֏yʲ-s��ӊ^\:h��'��r����T�lM�Q��3L�~���'Z6M!����yT �
!�B�(=�'�2d��&E&x�@ ���(,B��
�'Y�MCj.	�CK�/�@y�'��"�dٸ�xh
�Hґ_��R�'E�y�t��W�(�Qɏ�a��t�']����d	o�^Q����(Y����'M�p��� �~� �R��a��'������
?ل{�3YqzE��'���@�&vo��B�C�5mQ8A��'/b-�"��D�1Q�L
�a��Th�'�
e%M8Mo@�Q�GC�	-�K	�'�X�8.H�j <`3�"7&�-k�'��$���&��8����(D�qK
�'-:Q����3���"+Y5t�.j�'�������.Y� 7,X�k�L�*��� �H��+JQ�%!��X�ʀ1�"O��kv�,0
i8�)�n�<k�"O��j��
� ^� ��V�@���ض"O�Щt�"������4�\���"O� �@�.�����	@���d"O� �Aɔ��$=s���>��b"O^���l�B�ZAH����v�H��F"O���e�:1�( z�i<L��0W"O��V�R:�J���)�z��|z�"O���	�'.4�鲇P��d�[3"Oz�i�E�k�h���*��SF�!�D�֛�Pz��,���|��f8Ɇ�z�͍�9����/3 ¤�%���O� æ���I��]��m�3�R$V��m��Q� �����o���S�O�:��g�֨�쵉 �h	 ���~�h�b��c�ҧ�����	�;1��Z�a:Z��	P��^p�Ա*�>�U�EQ)TS �s�C.k�Ԅ�Մ5Z��\�h���sӐ �ܯE^"i��lXP�؀�xR*��a��O��\MBf ��IkHxش��FL�I�X�HRS�#��|Ҍ{�d�J�������3:>(���֬�?��k�����-Y�?1��0��)�%Hŝ���y�(ς+���8}�J�?��S2_�8���9>>�(ѕ��S��p)�U����d�Ob�����|:��?�"�s�A�9���L�%B���V��a��}�]*��:�u���ghG<N,<�;#��$Olrt�G'�
x�t�����?33�M�Զ�0|B�ዞ[���?L
L�;���	 >�\�{Ѵi �m{��)�(�KC�|,�lB�%X�udЕ���>iGsӀ1RW&)a�a����{��d ��ΓLj=h����y2j�|�q��	-�r��|����%��<s�A�*� za����$�4U1 $�>E��
s�՚�	�%P�����H��y"'-y��㟢}ڰ&�-u�&�T.�H.��a&���!���9�S�O!X�Qn��sq(D����g�0a�5&��(�yW�Qr�/��@ua�1M&��>�ulS�����O,��UB�� o&��V' �P:G�xB���O��pMXЧ�/�~��ŏZWV�9[�����'�lI��V�ul��Q��R�r�N�S�'�h�U	ǯ�L1�G�eg�H��'\r �Z����jR?Z�,�	�'x�e�0�� Rh�@r�֝R�Qp�'|����q�bD�V�XQ��'���@�زo@$!d� �b�d��'�8��L�h0Ɉ�)a��H��'Į99��� �>p�p�0 R�H�'Xd
�;�b�`�O[�M��'�C��!G#�ifG�P�~�R�'p���CQd��L�OK�-�'�0 �%��
�ʬ۴�	�F`����'���aQ�J��A�A��nC���'eF���k_�����AG�*P��=��':�P�BD��P��s��|��'����ށ �TY��/��y">���'���Y@ȠM�}�2a�!�DA@�'���s�g0�,�aa܀E �	�'9H F��֢�*d�9����'m�т�����w���GHH��yrJ��5jCʑ6$0��GȊ>�y2�ů	�p(�����E��Y#J���y�b�e}�vk�'0��P�5"�2�y�J�v2\�f��ug�)�����yB�ۨ Q�B\�j��ؐ���yb`�7܉�f� _�b4�e.��y��l���peŮFqJ��j�:�y":E��:$ƏH�X��Z'�y��O�c�`}��OAf(We��y��	"�h]+#䅫ܢ���h�R�<Q�)(i��i��6RL��xCd�<� P��ţJ4n\4�0̢ ���"O�I`�J`���)B|�\�Q�"OV�B��J8P�$=9D@P����"O��r���n�3�!;Y��4"O�\z��ݠ4��1ʐ����`"O������7Fh ��G�M-����"Op�۠�!4��	�F��D����"O��� l2L���CEE'���"Od����C�cv��QN�m=b�" "O�m�&Dq0�%�D(��+��IB"Od|�p�3;q,X�X

$�R�"OxA�+��F���k��(��ȁ"O��#�ˊ�`����!!�h��"O���Q��{k��ے�x��i+"O�ٕ!λ`�2 ȗq�@ErC"O�H�7(5Zܘ�%�	���q0"O&�bUhH��tx3�@}9�HK"O|c�h���ʓB�7'���r"O�y�#`�3,e�Q��Q�"$IG"O����o�w{ZP��Z�Vl��"Ol1�d,�
�8b�P<�Н��"Ob�r��
�Q	���p�xI��"O���5���J �	ڷgژ]v*��v"OqB�M�)c�C0^��� D"OZ���,�?Y��uG�ƻHj^|�6"O`�ӎB�Z!T	���\;I���C "O��]3tgŔ"#��v"OĜ�W��~�Z0L�-7}�q�"O����4i���O�p9�4"O☈�`��0n��H�L��ܒ�"O&�A��{�d��v��r	:��"O����mҩF��!Ʃ�4,��I�6"O�<A���CH����ovrp��"O&�34g\�Z�pLZtiI� ���3B"O�=
 H\�m�Z�:Ӈ0i�4�#e"O���QeP5d��%HV�ԅ��d�e"Oh�.ϭ�r��T��*�,x��"OPQ���	�t�0��K)Uu0���"OHp�ug";�-����,��q�"O��c"�("=P| �
��p�"Oؽ�ƨ%4�]���^�K�R��"O���(P���T:gL�"O��#�3/Ȥ���@O'L�~�BB"O�a�ۃ�N��쓛H���"O����b�<E� ���``�"O<<�cO� @z��kcK�-k�H�p"O�J2��$�X�9B��1�A�"Oް±L�&p1���:0z](�"O X3ƌ�:��`Е�֝(1 !�"O���Ճ@z*�����f'Z-X�"O,���Eq�<��ɼ(�a�"O�{�eB�o_�����T�=t>�"OցA��0%���1Ѳ�2E"OLhH�o�|w�h�d�����"O��1풠9���������cT"O��zS��y��X��N]�Z~�k�"O*M*ϑ�ۚ�;dLZÒ`�"O];d�A�C��1�.[�)�5"Ot(�&
��{F�
b��Yɗ"OVE8b�S�[$=�bJ��2z ��"O���u�F�]Q�����B�ys&= �"O 0�/���t������P*WHB�I�c5#u�R�c� 1pa�L�{��C�	�(9J�+=B��ce :b(�B�)� (��3�Ӵ	$H����"Oވ�t�&*�q���,B~��W"O�T[ oڼ"I���GIG3�u
�"O�4Z��`Ȩ�[�癅c Tӣ"O^Mi�Ǘ�)� �+�&4>����@"O�\�Q��9E��=#�`��|ר��Q"OiBaO�nߞ$yfo�������"O���\?<'�i2�hߕ
�L�Cu"O��+Y���QM�~�<r�"O��0EҖ4�",����1}���7"O�0�!�qt��a�&^���"O6u�sO�

��u�ޔJ�1R�"OPMx�-K�(3�ř� �]��iCf"O��s$��Z�ȝ�f��g.��"O���ùV�T�IԌ �I�87"O���q(�#	1p`�u钃=:���0"Op��+��QR�8��A�B)��Zf"O��CҨ�g���D2P�I0"OBAs"G�]oHU��-�%
��p�"O�|��⟉9�u��
Ƈ7�XA�B"O|�xe�ϖ(��
�c�ar�"O��ZФk�x�� -޴9D"O�yJ��-(7p@��frҙ8B"OB�P2�	�J��1!˶cp|0��"O�}�po I���3-�3^`��y�/�Lf6��Q���3��t����;�yB��FWr�da�8(kR�ju����y��T�@���6$����*�EM��y�K�p��RT��ga��yHӖF����6n-�reP�a��y�$�<��1��=~���A�y��؍\���X��
z���`s�
��y«��(P�U��o|^\�w��y"o�>}�� c#�&`f|P���0�y�BɵOO����ь'?.$K�j�<�yB
�,Ơ8�ݢ �2uM@�y¬S CE���"��Xv�Jt�»�y��Y�.�[�A��
����@LN��yB�R�,J�c߬}�2�R@�?�y�� 3�!�!o��0�#D9�y"BĹ|_�A�"$�4Y�D{����yBBI�-m�eP��'Q2}��.P��y�_�	�k�Fj��& N��y"B(:r�q�D�>f]��)��y�k�&JL��RJ>���c�-��y2&�#�V���C�#J�|�q����y��  0����D����h���yRn�?��!d�*Qj��J�yB�9]~����@5H�T@�Ņ�y2&�&�8��G��B�R5��<�y�%�T�Le��� <��9SA�)�y�!Bu�0�U-�%*�d�i�����yb@�	WC��@Ԣ�(K��BÍ�>�y"D,ir�"E#� ��B�K�y"
|5��)+[�jE�'&��y� �D�X*`�͘=���UG	�y2.D�]����/.e 2�E�H�yZ�X�	�DԞ_8��+ìH/E��y�ȓOߒ��̔7S�8���I�=1���ȓl_��rU+�8!���
d�X�c/V(�ȓT	@Q!S��AN���U	<1A�T�ȓn�m���Jm����q��/����ȓS��w�H":e���D&,�����&����A�W�D�ذ/߽"TBȆ�S�? .�k*(� �S�(ʜx�l;t"OM(:�h�(Q�:.\�x)&"O4��+��0#�D����eM{�<���L���{Fm��}�5�`�~�<y����BM�Tgة=ց@%A�x�<��߭d�������k᎜ꠦ\~�<�P/@\�{A��?��t�s�y�<�1��x�T�8�.6"�0��_y�<�c'7�F����@5{�j��_�<���ɌsB0b#��`Ll)t�E]�<q/Ƭ-�xL�3�UD���8Ѫ�R�<i��%4����"fNhj�����N�<� K�$�H��Fߜr� 7��L�<i`%͕Z� ��ƅ#��|�G��^�<9��
�#ֈ�(���F���E�]�<��!�j��98�%Y�f��%i���^�<Y� �**Y&��5*J�ة��KE�<��	
8]��)b�1�x x5�A�<�Ǡ��-��y �7�p�%��w�<��(Ǆ� ��Ƣ�5"�]u�q�<a$!ܩ΢��4F�pg�H�<��_�DĒL
c�ї1Dd9A`K�<���� Š �"DD��xӒa�`�<�g&�*O�|�dh�p��V[�<)儋_@�y(� C�<�r4��|�<��W,�³Ժ.RP�4�u�<!��+
Fp���R�^U夀q�<1C@��c��U��H´b��]���o�<�fU�Q	d$��f̰&��X�%�`�<���""�Je���,F����D�W�<�g-R�'z�AE��?20^e# J	I�<����Nʦm�6�:IK2M{���l�<i3N�<��)�_�\����u�-T�\뤭֒"�l��0�Z�r��!�%�7D����)�PlD��j��*|x'6D�h�#GF(*�y+�◬3�4�I �)D����P����6�ִwD�{��&D�d�C�K�Rl��EU�f�.m�1�$D�,�`���sߌ���NƤj��g#D�����
1�L�}��у�"D�d��$   ��   E    �  �  M+  �6  |B  AN  QX  �`  �l  �w  �}  @�  ��  ܐ  �  _�  ��  �  ,�  r�  ��  ��  >�  ��  ��  	�  ��  ��  7�  I�  � �	 n � �" �) 0 M6 g8  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�ou�!Dy�'�:� Ή�B�\O�|�����<a��$�+q��@rsI�E�f�W�]�1O���$���R�W����FޜO��'*(#=�O��)1�h�Z��K�`)����:o�.�<�J����<4���y`���`KR5��O��Dzr��`S��o[X�JC �+�lԛ�#D���5�^;Ki�e:	�L�� 3 �6D��@C�>y��HRc)ȓD�* �$?Oz��L�r�:M�\�H�| ���� d.���'�.���Ǒ����r�Hp*QGz�~RQ$X�E L��]O	�fe�y�<Y'�J�oW��`2m�V$��s��Any��'**��%�T�ncL�@���h���'���!#kB�踬�@ˊ	�2�#�O��G{��4F�R��F�|�Sm]�y2��6u��	��݆i����y��K�eb�#�-�b���q�����Otepa����+TJ y  �0��rL�C�I�t�@m��'[2H�U�LQ�!>Bʓܑ��|Zjͪ<\���,B�~�!�a�B�<��F��@��4�S�{hh����u}BX���ڴ��'4��'o��e�f��;i�(1b�蛞09����Z��� ��x	�aqP&�3^i^�Gz�D(O�e(P���0�2m����
ba���"O�mkF��f�-[����gX~��"O�Q��gX=L�(��kL�*mA���[ԟ�?E���P��,A��ޛg9(\���C�̄ȓy���C&�6��[�M:_�,T�ȓJ����X�%;4�҄�B�kTL���	|�$�8v��Y��l:n�뀣�;RV!�$ ֒��O]�6ě� �HT��\E{��� �QZ'���Ԍ����<	���"O,,�p"T]q������^`"OL�:���\�Pq��@Y)u��x�&"O�m�S�O)t�~T�%IM)n�-J�"O@|�㢇s���ʡ'K8IO�ܸS�'b�O�l
&C��~"��ᐙ;�fY���	4$E������}��p�'l���L���<}Bd!##,h@���W^`򣉒�yRN�C�y� ��"P��)��
�y��	�c�e�хI�J�Y��y���QĨ�J��43�e�ъ�=��O��~�ѩ0�IBա���@�@�P�<0�C!��8Ӵ!�0r��ЀRD�q��D{2&�r�P�;��O�_^�Qv�@��y Y,a�Lh�ؠden\����yB�U�2�C�iX`X������x�iNx�(Q�ԪP�1�C`@�p5��>y�'�R}��j�Kn�0@��G��%KÓ�ē5�����~YI��������d;6�}��!PdsI�b��E�3�\.I�����hO�>�1	 �p����ʚ��N�x�a2D�Z%mA<���Ec�u���c ���E{���\�d<:��$�%qp�y� ��!�\~�R'J��JT�cԦ<!��Rdbm��FC�^A(���B�!�D� &��59���XO"���A�)8!�� �Z�� �Q�8� �O)!�$��V���ʡG�=,��cOE�	!�$U�"�Z�!�A� y(B��m�+�'a|��V��mX��	� ��Qa�R4�0?�-O��ST�,��88�8H�
��"OZJ3su��sU�V�t�g��0$�,2ٴ�M�۴�Of�U2e�ԑ+!ƅQ�)B���'R��PK�0wxfK�"��m�H��1�4�MS�y��D�ȟVD��k�dU @�e�F���O��~·�8~X"8�aÆ.VJ�ڥH@y"�'���c&��*`�!��	x+̪>)L��(��Y��i�J&�9���~m
GN:D��C���"t���ԩ�'p����e2�I�~�O��˂?2p�`"�_T���' $��`�8x
,�S,��jl�<޴��'꠨�㉁��(	�N�(��l�eWSdC��#e٬][�N�h~�h��U�B䉷A�l��e�zVLaei�n��⟜�鉰n��A�x2THU&^�X�B�&7,`T�w�l�J�y��ij�'�M)tΉ5r�a�7�M61Dp�'�(�I�X�91�ɑ7��),H>�[�'%bаf�� �.��vK�:��p��OƢ=E��&�:Kw
ϝ]�
 �3*D��yr�ΆZ�>�wO�Y�9�ee���'m�zbiW�8\P��B�W@\L��/�y��R�*��
�2zB�t���7��*�S�Oav���?$8��B Ts�@�'&������:������/:����y��'��XB�EiRm��K��]o��
�'6��*�,X�� P`B��T���'Ax�oM�| �ɶ�A�TA4���d.�n�;p��$ܼ�;�KDu��Qi�"Ox���S��ϟ,.�~ez��b8��C ��-w���Gt�<Y��8D���Q�5$[�x��h��W�)D�(����V:��j����T�lK�):D��i���>������[bt@��B7D�� �t)�ȍ�F�!/S�D3���"O��mʀ*bfu����4j.��(%D� �pI78�ޅ1��t�cm&D�ȳ��O�>�z5ʀJŘXSF� �d%��ȟ����_�)7(E�KM�b�S!�x�'D��pN�:㞁��f�$%�j5�
���d�L����FL�D� x��T�!�$ƦC�&qb��@�(:�V�� �!�Dߋ{����6<��E<�!�ĉ�^�z���eN� N`��7�"f򜔆�@y@�� .�&u��|iv΂�.�,|��ȟ��OH���� beHT�dO��*t�ҝI��	��.�~�'���l��� �D�#s���'��l��] 5����╀e�Bh��4�~��'�����$ {�̍a�_��(�K���4&��?���MBx��˖� sbi�d++D�d����84�e[W�J6.���%j��O���ħ��/�v�Y圻��K�*��hƜB�	]袍cV��;����5�Z	dc��$�x#�'�ayb�����Fc��
V���w U���x2�ޟ.�H�3�E�Z���� �3x7(6mh�
���E�8��5��ǎ%nؾD2V,
�T��O*4���	A�uW�I2��:f��P k�j�!�ǕV�����F4$����I�!R��	�HOQ>��m���J�{lA�;���,5!� T���1��i�ܠ�M�*P4���>)'*B;F0ѡ�$�p�ڈ'�F�<�LU�Z_�H%	e��c���x�<��ϋ�I$t��cO�Kw|Yc�J�O�'1�O䠖O�h�O��j���X����h�)+	�'���A��"�b���*^�T�"Q0�Of����>�Ģ�f�!E4����֠i!�3C]pQX�N W>�i��a
�QP�_�l&��g�3�Ha�O���%:��тact�ȓ*$�(+t@2*K>�9�dܨa���ȓ5ю��@�4	�2�I��	�=�(i��c�����"���&���f�$�BI��%s����*Q�x�K���"5�^Q��:��Eɂ��0zGv�TK %�<��#f�i���
��TeM�kθ�ȓv� k�e�EB�䢔՘C�jy��)V����H�pE<-@�J�B�e��I�v� ƣ�
�=�b�8�Ʉȓ/�<ٙUn�
���u�K�XO�ȓd�S�+�{�	�c�%z��p�����e��Y��9&
�t]�I��P�� 1�(Y��Q���A?� �ȓ-��1Cdk��Z^�5�7�2u��Q�`=��NX$!#�$�&mC��Їȓ["4<����zO���&���M��V��U+S�0/bU@҃<7��p�ȓZG�ي&�^?�|��6>g���z<l	�V��$�Z �88Zh�ȓOS��r,ہf�ԣ1.�2fW�Ȇȓ.��-)��C�c�$8R�iäs"`}�ȓf�&<�b�
.^���c��%Jm���ȓ5�ڸ	g���K�����ʉ"6�P��ȓ5���GF�e��}����&Qv`L��:5�h+A��:��s���W{����qr0�Q@%yp-�P��o�&��ȓk�y#Re��.�ܬ`bG�5}�����}��)#ӡ� )E@�0��I�Go����\V�0Ň�e�Nܰ7dF�kԵ��%�܉����2�A䨂-&� ���S�? �Hg'��Jd ���3�=�G"O�a�#��//h��Rl�Y(܀�"ONbC�$�U�jN�J�kw"O����KP
M�`)$�Y;�"O�Qq�ʜ}P���g�T�ju�6�'�2�'Gr�'m"�'�r�'��'�048�̂#g�h�85
W�0>�d���'�"�'���'���'%��'��'r��g�<J���u��7�'>r�''��'���'���'�B�'�1eBϲ	;Z�jFk��(uڃ�'.R�'�R�'*��'��'�B�'a�a�T�I8*hⱺ&��4=�p�1�'�R�'$2�'�R�'}�'8r�'��Źw�P�mx"��Y�Lˢ�'��'w"�'/R�'ER�'�b�'���G�	S �]���+n�� #�'S��'>��'���'���'�R�'bP����F�n�fc7(�i���'l��'R��'���'2�'�"�'@���f��A�z��1� ���`�'_b�'�r�'�b�'���'���'"r�:�eć5����"xEC��'V�'R�'jB�'�R�'2�'���$e9
��	X���?.;r�Y&�'m��'���'���'���'1��'cB��.�t��1qs�ԧ%?����'�Z���':��'���'�R�'u��I�,t�+���b����ETjt�'s��'X2�'�'>�6��Oj�DX
)��X�B�?*"ts��
V��'��]�b>�7�Ɗ�,"NlD15%KMZ�P)LD*��2�ONlp��|��?�!
�7J Xt�U�O� L`����<�?	��`U��ߴ���q>������� R�Q�͘t�n��@ I�1#�c���	KyB�`�v�8B��I��@�6��37�QQܴGܴ�<���$�f��n������.[�#�P�����54���$�O��	_}����H��<O�4R����ZH��S틇d¸D7O���?AF ,��|:��-��A�PĎ�i.BES�E�;l�Dp͓��d!�$�æ�s�k:��8]ʦO�5n�̉��$7X]���?	%^�\���������3#�vD"�m��"?�i7f��3�����$R�b�<f�c>%Z��'g��ɮ!��LCTG$�XD�cV�^"�'5�	՟"~ΓS��Š��_�����)&Ht�rF�����D�����?�']�L9���ނE^�%�&���#��}��?Y��?�����M��O��3�:倜�7 �G'�! Mn�6.�(rVʓOl��|����?���?��t��]Cu�͈P�\��C�A=.�dQ�/O��o��J��u�	�����j�s�$@����fS�0;Ei�+
�ap�����	�kڴ
M�����O���ـBO�	2�P{�,y��	�(��ʣ�J
U���W�� j񡌭<�뎂D�	�򤙇)\ȝ���s�E)HM�Isa|"kcӴ�Jp��O���PB�g��h���%kHh�3��OmZ]�1�I��M#��i�\6 �>ݒa�Μ)n"�aj$O�L���v��D�O�P@���J׎�<�'��;\8#nڠ�ע�*g�n�����<9
�Fk� \�>`3�C�����?����v`A����즩$��a3��z\�YAI��3����CZ���i>��vȆ�n�5l�]��00�tH�Y�j�ekf���X�x�	p�Imy�I�lyK���ڪq&��%~.���4<e�Ě��?�����A�UoQ:�c�m�j$P�	��g��'���O�D1�4�~��2EZ��bC�{��Y���5�N� QoR6���m�<1�'x5���t�r�R�겠�,[����0��DU�������ݟ��i>�EO˔$,>��'^7M
X�Q��e�)��)f��E��� !�O���[ڦ���Py�'|���?1��͌=t2V \��a�3b�0T�(�d�O,��6I�=v���O��ɲC ��4_�<" ��q��a0Q(k�Bh�vHt���'���'�R�'�r�'�S2=dL��`��'����38=�ٴX�rԉ��<���%.I�?��4��w��y�׫H�!�zi�S���Wo�aC#�'�B�|�O���'LB�AǮ��y�>wB�%���E�2��X�ᆙ��y2$[�8Y^����?�s�@�<�*OL�D��>�Y�%�#���$�Џ �N���F�O����O
 �F�<aD�i	�Y�G��y�'��D�2(��p#��]H\8��|r�'������C�:8���[�,͔g�����48�ퟜyF/6{<-"A#9?1�'i�~����P�t���&��J+�"h�c�7D��ZPfM(>P������%T����쟰�ٴn��a���?	��i��O�n�0Q�0�2C*�;~�V zs/C!
���玲pߴ6��f�U�]1����'1�BQ�{M�өp���Ŧ�;>�PLz���+	]�ę|�V�t�IПd��џ@�	�H�ɓx�����;�z�⦌�sy�{�&�i�cʈ+����O:������D�O���P�ǷG򰚢fP�),�ɱ q}��'C�O�	�O��d�|�ӄ�F�[���:��{���O�\˓X�D�FN�O45;O>�.O��g#�.0G���"�I"S�: ȳ�'	�7�������05�6,�螳��i����bl�DM����?��X���	ߟ���Ѫ5#Q�#�0�r�씲J������3Z3��	矸���	����<y�'��� P�J�k��"����6�1?+
�j;OT��䘖n)�X ��B8fyָ�Bh��7���$�O6�$ɦ�R�a?R3�i-�'��)٠��aDly����9;`��6�|��'���'��X&��y��'��)�P��f�l��H�5l���_���������d4�	�ga2�I�*��8�2s�4Q��#<���iL���t�'��'��S�	�T���Q�`@vǆ\.��.^����MK$�i�O�)���0�ѧ�Z.�<��/2�A��U}R���E��>����1��O�48M>���v;vP!d�L�
'����D�p<�4�iy�X�Ǡ� -.`a��aͼ�x!�$�)z	��'lr6#�I���$�O�`�(�
RrT�Y�fW	�����O��dO�A;��@�8O,�D�
rr|�y�ON�	E�V�94���}ɚ��d��u9O���?Y���?����?1���ٜ0������4�]K��ͣ��lZ>X�������?���П �	��M�;pEn�(ƻ��aKůzP���R���?)��O���'8r�冘9�y"�Cl����I�W�TpKvc��y҆_2X��E�I�d~�'���_yR%ʍG�(�bҠM�@�$�����0<i�i=ڤ+D�'i��'$�Kg��/{²t
ӣӏU���e�D�l}b�'��|BO:�a"G��$�l1r�d��yr�' ��@�]%Q2��8�W����v����O�|����1�xa�a$ט&>�a��"OLyQ�ʛl��hS�[{;����J�O&ql�bt�	џlc�4���y�O��m͂h�EG��-��/Y��y�h��mm��M�$�7@d8Γ�?1�.Jp�t���6���Ya*�6]*j���D�L��A�,Ԁ��F"_]<�+O��p�����pp��F�X��{�� sP]�Q�a�Q���Y7b���ں"Q��yEiLO�©z��U?��K�Ǟ�M��d����M2%#p�ݴ &�i�	�;6����rژ�� �b��7�~��Ӯ�#�����+8���kҲ$����ߒ�K�
����K��B�b����S�`�|{�)P�^�,��G�ˠj1E�f�˰	�*uIEM��n���
W�V�t:��;+W�B�\���G �RŐ#j�|d�y�cCV%B��`�Ѫ:�����~�\��OX�������'�Ik���&5V���ןq-"�{޴����1��b?�HSE�0p�x�چmU����%!mӞ�U���9�	�D���?��M<���9j0�S#	�����ac�K����i[���֟d�tl�,&n��3V�Ӷ}��D�"���MC���?���6����x��'���O�Z�F�G�uز��y��DO(_�1O����OV�DɣD	�1�7 �^lȽGgȦL�BTn������-���?i������%ƿr�6�(�,�5���%��d}B!E���'r�'%�]�4gH(YEشk���ae�}��dȀK採�M<����?AJ>�*O� +�&�-%:�i�M�)�6�je\�"1O���O����<9��\�6��A":�������Ji���I�'�R�|2Y�(1W�>��L�*�J� s`E�z�l5iSE]}��'��'��I>B	3O|�F�����H2��R��:���v����'iBZ���')N�˟�	� 0�3"^:B�u"��&�7��Oh���<)W� d��OZ��O 0��'��$�p<PA�Վ	�k%9�<�B��K���	D�E�F\q��QNE��P�H�K؛�X������Ms�]?��	�?q��O��c�O�A%�=P����:�:=�V�iz�Ɇk��"<��'Of�0��_����#�Mb�.qs�iѦY�I�p���?�9�}2�-<Ē� �O�.�p����,=k�7-�)�"|J��xI�IkLJ-$	�4kS��.^6m�s�iU��'o��3O��O���O4�I��T�+b]�9�6���l���}�F)��'���'xr�K�hl\��%ˆpΖ��w��6m�OixB� r�Iڟ,��I�i����d�#D�e㕭֥T��iH���>٥kf��?���?��?�ߤn�fa��i�12�L�a�Ժ;�xÆX����̟��	f�̟��I�	��,
�)ڙ_�(�I�'F��2�f\��?����?1��?I�������2��I�G0D!R����M���?	���䓣?�M���%�Ȧ�86�G�O�Z�"hO�$x�`36�>���?q��?����,E���?9��[>��bE�Zd�.�:�k�&mM�t��i���|��'��	� D�O��N�����%-I�1Q�L�վi��'�"�'S�i�'��'`r�O�^�E]�j�pqA݇X��i0�(��O�QT�DxZw�x�90�I�<�^iJ6�g�
ߴ��Ĕ�_�����O���OT�	�<�1+�$������He&��%�
Q�>�o���I�L}���?�~�@�Ƚ-{.Q��1Z���[ JE���w�O�(��ޟ����?)�'~��'w�����B�w���E�̚�u�VX��(�)�'�?­0̭����P��q!�V�@D�6�'�B�'�J��$Z���	蟌��`?�b&�Z�q�B �5@p�[���ͦ�&�(���ޱ��'�?a��?A��I�G��Lb �)4����P�<���'��a�T�������Z�i�iYc�ł�2�p���z���h�>�@�L����?���?a(O������*t�ȑ�7����n?@��˓�?���?�O>����?9t�<�,�gH{\�u���i�M�����D�O*���O��[0���π F)Wg��x뀇 %9�r�k��i��'�"�|�'���fJ�DZ�8r4D�Ĩ��e;�m1�	� v������Iܟ��'�E�\>��	9yIC�׶9�$���^�x�bj޴�?�O>��?	���6��'��hi'�^g��;G���~ɘݴ�?	����-RG��'�?����ӎH#X�i�MG$w�4��u`��5�'���'ZU�5�T?MCB�ӓ)�.9p�OY�D�	���c�*�`͊0:��?����?a�'��Ƥ�J2��(�b\y�j\�>�:��iH�'1�!������6�ѐ�
Z� ��֪Ȕ/���C����'���'���[�D��ןL��E_�x���h�7I�DQe �9�M;�ժ�������� e&���Dj�:w����e�Úmd�o�����ȫ������|���?1�|NvL�JU����	��]��V�'��Z�Tj���	�8�I>'s���֬��1�Fᛷ��
U�u�ܴ�?��	�)����$�'ɧu�G�����C��>t�X��%���?*O��D�O�d�<ɷO�@��AI�|�,=j��i��Ș��x��'��'��	ڟH�I�� 3��?[���Z�'܏)�4�k�ĉ��L�'>r�'����H����O��3Ttr��(K@�1� �����̟��?���?���BK\l7_���Puk�+cQ��J`L�O��<9��-a��*���r����"��T�� �Z�l�B��?Q����U3�J|�	���  �0@,r,BB�T�B�D6-�O�ʓ�?������Oz����k��(Q� �����s���vI�2i�'�2�'kTA��ʕ������3��Ѡ�͇;P�H�C�2Rh��S�ds��µ�M��V?y�I�?���Ot(�*__�N�a"�C"^K�!���i��'U�!6�'y������|n��D?���PB<��|#���8]��6mZ� ���OF�d�O��i�<�O>�dXvO�vJx���/K6<�ƈhӦ1Xd
1O>5�I-����ЏԄpLՃhZ4zi\E2�4�?���?� ��<%�����'{��$m�<��,�1WU�z҉5^U>6M�O����O�1i(�G��O���O@y�V*U4Q�̽�`�W��|�C�	æ����(~f0I<ͧ�?q����U�Q���5C�.^�Ш�&J����o�џ|��͝џ������'�IП�Z��9y~���@��W�r%�Fy����' "�'�O��O��{��|d���F)�*y�R�q� ��t;���OX��?)�A������1I�$9۲+V�I@̘r�Ӹ�M����?��B�'��ė=]\��ڴ[F�c��7��y{&�����?A,O��$��'�?�sL[�o���bLƎ(u��Z�b� ?�F�$�O���4K\)��x�aB�6#���6-�j0{ �H�M���?�.O�)�c��[����s�Ѻ��*U&
a��Ǉ,H�6�"�c�z��?��orN������'��1?TV%�jXDu֕���+a�U�'�r���-)��'���'���R��ݴY-Du��V}�����(bLh6��Oz�D�h������-T	��'�#qV�)Ю��Fd+���'r�'��Y��T	����.�*"yV�X�P)�p@�iꔔ����☧���d�z�2���g03%���T��{�PlZ���ޟ ���ϧ���|
���?��M�0
���O�lȆ�0�� ����'Z��'KH����~Γ�?a���?1cԸ��|�f.N2��8`K�'��6�'>0D��H8�4�����O���,X��H�P��\�Wl02� <�»i��LM��T�H�	���	Ryr"Ԗ*rM2���C
b	ã�PA��N�>(O@�d�<���?	��A�"���Q����,�H�����<���?9���?�����Db�~��'j�<#�ĥq .�����Fi��lZ\yb�'�	ܟ���ݟ܀b�~D��P� �-�Q;,=1���Y�	П�����'�x���~J��p���S��A�ؑ[&1fh�M�Idy"�'�"�'�5{�'剦"����4�JY����W�fM�Xܴ�?�����D�$bl.L�O*��'^��ҍH� �*��	���E Y�jP���?����?Y�,y��O���e�!�� ��l�� T�_�6M�<Ӏ�R��v�'���'���%�>��:Z|5 q�3x� ��Z�z�yߴ�?��GHyΓ3��s�t�}2�+N��:-���e�"�
�!ͦ�cd�M����?���b�X�D�'I��[�nV�jbQ�DK� �i��q���*�6Of�O��?A���Y�Ny��na\�9���m�:��4�?���?1��Ap���'���'2��u����h�9�J��YhP����M�����e��?��Iן���d��0��'8Q��*W9'RRq��4�?��L� ��	ey"�'?�I�֘~5�ͩ�BВa��ܣ �q����h���?���?����?(O�����?$�-�EL~���
M�	�n��'����'���'�����}\����$�,�v�Зb��IJy"�'��'(��76�2�O�\�Q��� V�K��:t�l��ݴ���O���?���?@��<�1'����KE�4����4a��nߟ��IџX��ß��	YI�`rش�?9��:�~����3:��� �#P��x��iVr�'��U�\�	�� �=�BL|���ٕŏ�Hk"P3�͎�E������	ğ@��#���M���?������ �������G��\۷�4T��hqոi>W����T���]�i>7mM=X����3Cip���'*�n��`��7�O��D�O�������ЃS�d�k�@�52d�����EY�y�'k���S|��'�^>�L��V/[6��1{�L�/�p�8��i+���V�q�f���O����:8�'^剹z���rd_]�4d�+�0j��Y��4uR6\Γ�?.O��?��I)qzTpWH�sH�ACP�4m���ߴ�?	��?	!����'��'@��u��J�Y�|�
!�U�Yw�I��OO��M���?Q�.����S���'k��'�f	���?\��1e�X!Fƨ���`Ӱ��|�勸>�-O���<���BZ�:�V��P�X>�����lLe}�f�'�y"T����ן��Py�A˼9����r�����yS���N{*I��b�>9(O4�ħ<1��?���?�̘K�c�p��-xR�T*�k7h��</O"��O��d�<!I����Iߞi!�j�4Nr$�qb�$3�m�vy2�'H�����ܟ,�Lk�x��%l� ��� /D51��!�M���?)���?1,O��s�`�@���'a��Rv��bW�)�֠��y�lJ�j�L���<����?9��?�T���?��'�2 Q*E�k������⒪�%�M����?�/O�$��H�T�'?��O�F4B �d���*�������B%�>)��?A����"a�'���'b���D�^ ��L� ��,��lXy�EI�2�6��O����OJ��V}Zw`�`��NBm�h�Gn�S0���ش�?A��L����d�}:�O�i������?��D
L̦%�"��<�M��?	���ZpV��'D©�@�]�	;�L�1(Ȥ�Q�gӤ(��=O���?�����'� ��$앴],�
�ǉi���#Bd�����O���F�'|���']�I՟$�[z\H��ڑv�����]�p�'��	�ך��|���?���02�'*JK �91��("��*�i�^�<߀듶�$�O���?�1M�5�w���@]d쒐������'���'"�'�R�'
�s�<��_3`*���0St�)��(|����O���?1)O��D�O�����A��+��O�A٢Q
2&Wu�Yag>O���?���?�+O����M�|"��]@���P�]�`z<	U��X}"�'���|2�'��H�9:E��	Fq�}sQ��y�Z���'
��P��?���?a.O�cψk�ӝv��k�d�1py��@�M�v=��z�4�?�N>I���?�3��<9J��*�ď�c���'�F�<����ԉr�����O��r��՗���'���ŏ�&���W�q�@h�C�\W�O��D�O�mz 0OX�O�S������
��h(�'Ԁ]��6-�<Q��	 V���L�~������� �K�6d>ȋ֥�N'Z�g�o�z���ORY8T��Oh�O��]Cu��++*����ǝJ�dL�w�i�eQ�.e�,���O�����$�$���	�K�6 	�j���`r��@��u�ڴMWtY��	�Oڄ�%�_"@�
��	]��q�Ҧ��Iȟ���75t�KJ<1��?��'�-k�(�pK9@�� ���MkN>�1���<�O`�'�����k��f�D9{%����7�O4�qG�`쓽?�O>���J �Ӭ�5fb��G*z��'-0��'X�	ȟD�	ڟd�'Y.�(�ʻrk������8��rCn	0֮O ���O��O"���Oh,KW�S�?ۊ1�U�YcF��i�X:��d�<I��?a���B�E^�̧iFV�9bG��ȕ�f	�/:ژY�'pR�'p�'qB�'n����'-��o�[��K�Fą�d=:�˿>9���?�����]L�$>��"��*-D)�!O��u�*�#�Q"�MS����?Y��|(ʭ����I Qr��A�՘O+�u�����7��Ot�D�<�&��)Me�O��Ob�0g�//rT(�iW{���_O>���O���-�O�O� t�:��f�؋`�@��F��z0l6��<�f��$mi����~*���������ɃU�R0Z�͇e��� �b�<�d�O� �g��O@�O��>���ܪ{�e���Ä��i ��r��`����O����@$�h�I�2�s'�"I�r�#k޺R��-۴#<�QY���S�O��L�(�t�K��@�~V�͂Qk��Fd�6��O����O"Qz���]��՟��	c?!PeX������O��ڽ�p��ئ'� �#HP���'�?Q���?V�_���h#�ş�>�z���&N�#K���' >LZQh5�IПP&�֘�1�^��B/L�z�\p�5G�+�|�E���M>���?����:O�v�sĠ��c�r!�/�~��6c��!�O`�D*�d�Ob����d�4�Q�P�n�|��A�J�8��R?O˓�?A��?,O�����|b�CS�1J
�x���
��|K�e�J}r�'=��|b�'<KԊ �)Q�;0�0©O*?�^���֩0� ��?q��?q��?D�ٞ����'��[�8ڒ�t���·ЖU?*6�O����O�˓�?� �E�|���~��̈!P���T��c����(��M����?1��?1U�Ϙe@�V�'n��'
�4c�azU �������Jr@.@7�O���?�͘�|����4���!�� ���%��<����.�M{��?�'���6�'$r�'��d�O�M��a�dL0)����pc��'/t���?��
��?����?�(���O=X�U���/�Aj��#��5��4o��`���i���'�"�O����'���'�B� `����M���'�)<�E��i�6yP�'�ɧ�����'J�8+G�?���i�&8hOn<hdca���$�O��d�4��!l�ڟ��	ڟH������8~T�3�QEV��"
�F6M�OD���)����?���?h�����z�JsF�Y�;5~%�ưi�����b66��O@��O����A���O�Ъ�� =-$�@k��ľ_�N��P��zu�w���Iϟ��I�X�Iny�%ά\�+MХ�@@��_*1��Is���>!.O���<)���?���y�$��t�8+a V�_7N�(x���D�<����?I��?9���避9pqoZ�C�d(k�4�\Qr � �*�Qٴ�?����?���?.O��d��|��X�NP�]`���>+��4ȶ/[�x�l����������IOy� �Z�꧚?qwa���E��K�Wvh06�ǒj<�f�'/���P��ݟ)E�&?��u�2��7\����J=	J"�����'��]�`ä��&��I�O������t��լ8��pƀH4rT�ӣO^}��'E��'� Ī�'�rT���'*n��K�n��1�b�; ��8I�Z<nZyB��*��7m�O��D�O��I�x}ZwD� @��w��%	�L�dA�l�޴�?���t��X�����O�����˃C�*����R�Y�"Y��4!b�l�E�iB��'W��OG듨��Q�0Ur!�Ʈ��K)r�c���*���oG���<�'����d�ةs�Ϝ0,����U,U�:|�o��������G!�<��ļ<!���~E^4Z,E �o_�*B��A��ȶ�M�N>���<�O�B�'����x��0럘EI�١�D�-TD�7��O��+�({}�T����hy���5��+���� ��f�x����M���D� ϓ�?����?����?�*Of� Vk��;z�Q�!��3��q��/��S���'2�	� �'3��'����]������4���7?q܍1�'���'���'�"Z��c�kO���\:���`Μ7+:��fRc֖n�Py��'���П��I��<k��>I&�؅63V	K�M��O�`@Y�"�٦�I��	ܟ@�'��9�&��~��bvAT	B!����3�&������i�rQ�4�I����I�lz��~�ƀ8�`�Q�K׽I��\!ĭI��M����?�/O^QI0��\���'V2�O>������N��Ӣ�!R|��8�b�>!��?��0�����d�_c<n �R-��1P�!E��M�*O��c�LϦ���՟$�	�?q�O�.%c��r��Ȭ`T ��3�	�b�v�'��ȟ�y�|"�ɖ�oe�9����u6����)ͮ?�����"�6-�Oz���O
�	^}b[��+�	N9���r�k��ITΝ0�ML��<���?�����O���k����-HǤ9��$'��7��O����Of�9�$Cz}]�H��B?�S�+Q��R	�1���u)�ᦕ��wy�̉,�yʟ����Of�?������:y���P��u��4�?�&3���Uy�'u��՟�X�(��q	�D�;j|�xpE����@N���<a���?I���D]�}}t�����s�ukA`�,	|���GXQ}�\���Ity��'�R�'8�G/��w��у��/q����f� ����O����O`���<is��@8�)�q�^�P��K:���A䬈�^9��^���fy��'kB�'�.�'�Is�	��Gj��s�ěs�$l����>���?q����Ĕ�Hk@u�O#�	Ѻ/)��2PM�.M��P��i]�w~7�O���?����?����<���?�n�!~t�@�N�"�3�N73����'Z�Y�Lr O�9����O����<Dȕ-_C�*��%�sY�%�T�S}B�'(��'E\�'��s���'ɬh�d��<\&��e�3K��,m�Uy�B.��7��O����O�i�s}Zw4�"cgՠo4�X5ᄨMf�9{ٴ�?�c	D�'��IK�'z���Ђ�[6��B+Ax��mZ�M�I0�����Spy�P>q�Q�Z<�`$rb,Kg�lL�����N���b>��<Ql�`iݖ���qu�._�ژ��4�?����?��nO����D�'�����,��J�"�# H�3Q/�A��c��{` <�I؟�	�
��&Ra��K��\��M��;��A,O��O��|Z��6�B�QC6�
V��({A�Ƞ5�Dۊ.	�	̟,�	�� �'7�% �+��P�RB��%����D�c�x�I՟�'�=OhiB4�_K	.��3�);��b�W��'���'-�/$�����/Á{,�(ҫ�u���Ɖ�Jt{7�� %<���!d!�E��&�� ���V$D�;��"�qO�V��/��i�
�㝔d� �7�[��p(c V"5�j9��LV�p�,�!N�8XU�S*��`ݼ�jDL�1*��i�[8њ�kKY�L��m/4$��PfȃR�΁R�̋3��֟%w�$��!��}��)��c�>�@�e`��n�u��ԤC* �`I�����	�w�}{!�j�He)��")����(!�5�0��`I�@m�EC"�݈]��i�|���
)|����"��Q��8]`l�O�hp�,�(Ȉ���ZR�nZ��u7��Y�OI4��UbάvX�Y��d���M�X����O��d/ڧ�?9f�B;7P����V:pTيp*g�<���Ĵ����,X�K����d�h+����:&D��1���s(������mo�ȟ������[?Ĥ� ��'�' �w�v$�Ƣ�Wt��L�q��H�lG�HM���'�=�禉Ә���2���o��>�\"�D"3���.�-�������5�3�� ��Q;z_��@)�1J��@�e
�O����O��D�Oq��	<�D)���ٸ3�N� �ĩc�@�Vh<�4m[_��)��L�KC<�"Շ�y~�$&����<��g�x�MYB@��_�ar��ųǠ��gQ�?���?9�x���O���z>�!!��ۥGNx�����Z�d�C�	0��0��� j�r��N&_�p��!�4�ե�� rńH�42x H%�� NN����O����OV����Ȅ(���K�>9Tx����$K!�2�|����\!9 �\�hQ9j�1OB��'��I�@��B�O��d���� 2O%}V,��iT�@��d�O!*@A�Of��|>�Yq�ܹ54���M�
p�=o��z����FV?{7Di�ϋ�`-���� c�2eT϶	c^1�Gr�R@{4��t�L��k��M��d��'9�]
���?y+OJm��$�pG�m�%m�%v�H�{��5|OT�S��V2V�h�X�bR�ckʽ9TO�MlZ�W?N��C ���0��ե"�"�	}y� �s����?Q*�f�5)�O6(�����1�G�sn�ܓh�O@��vZ�(H�DB$9�ܬ�p�I˟ʧ��I��_���!��L2!���(��+o�Lg��	b��?&wN|{6����H�<�a �#��A�Q�6]!G�>)7�B럤�	k�O�rǐ�f��֨u�*����y�OבlQ9��2)q�+��0<q��	�,qn�k4��`88�bʇ9H��u�ڴ�?����?��U9TF�
���?q��?�;%Y���ZR���ԕ*��)��y2L�L��I�=l��Qv�Ÿw����Ձ���YӌM�G�ax2��6�(5�4(E�+�l�.J�B���24L�Oq���'���A&&24��,Ѿ�h���мGz���	�9��I7�V�1t��(_z���HO��oy�'9��2�Ʉ��)b�/� 9, �j �J?rd2�'���'��ڟ8�	�|M�m�p+6c�:�T�!U��@QҤ���>�PBT���,��S�`/=@*8
�d�Q'Ȝ�1��``i��I�Q'��t��60�� �D0%D `C�Or��O��D�<Q���'�q˷ʚ�)���;��ȑ�bi��'pf��ש�#j�^��AN�sO���y⮱>�/Oa0c��9�	ȟ��#�B�q��pbH���E\ʟ��I�Lk��	ߟ$�'Xx��&�'h.a�c���,���܆xl�x"" �4E��*�%<OD5H�.� x���$��Jض] ���-�Nl	�!�(?��ҁD��p<1�%ןT�������oX&�C���kn�А�s��'?"��/cƼ����� )�QkVLߠ=�jC�ɐ�Mc6�N�2-��f�>N���<Y/O�#�^d}��'��S�F�6q��?����w���lR�,`�j�	���Iğ�H�#��!Ŗ!�����I�d�C^6�$r��I��L�3�(8��[�@'xLHצ����	"3��L�L�Q2�)�v��7d:�j�̔?��S�� ``�((o@�w꜄�2�'W؀��?y��i�OvTa�f]Lw� %�F�P�JI��"O��H�M�X�R�s��B�"	ǓIj����D��"K���5;�:��)��$�O��d�0ag�l�gi�O
���O6�4�`I9bK9#������ jx���`��3��Rq/���D��A�bc>�O~�i(�x~ ���F2o�<�A��F����t���hz� �dq��'��Ђ�OD%�1�mעzR��'�B�'�t)���������O~��6⌚O�[&��9�θHGE"4�0����j���sƸ�A�%?a"�h�U��-�O��]�V��X1D1��o�("��p�֟p�Iޟ��ɏ��)�O2擀;�Ԑ6+=/��UP��	��(d��T���mT@%��0�n0iP�9��
3���DDSS�����I���<	�004�� �	��� ��6����x�I��H�'�2�d�LC����gt�����2 ۘ���'v�}��AA��h�Ń� �yr�>	(O�܉�������՟�-�1JOp-
��ؒjy0�� L�ʟ\�ɧ4������,�'h.��c`�X�YY�8��O"<�'ɀPM:52BݝBuKa�'G��Ї��C�-6��4�0��< ����>g�y���0O\�0�'�"�'򦟭N����F�,�AH �2nk������?E�d�N!	@��brLY�9%�0��o��x�lq�(f&>K�2�H�e�y�ڇ7O��H�R8 �ir�' �,^�d���?�|գ�m��O\D��lC�O��]�I��"X5����GI�<���S�_>A�� g�PeP%���sr�p��8}��؅V�.p�N�Z��$����^a'��}��x���ƴ`�Lӧ�'Mӟ4�	C�G�3� ���LM�A�@`��J���G�$�O���Dތ,�P��RC�3�`�G��axr�;�;�H�;Q-AR���0Ȗ�n�<Փs�i$B�'E"�7y�����'�"�'��wB��H�	Tn��h��2cf�$�c�3��_�$,��m(�3�DU
!��)�.�-�TJ���h��% �k3?���Q�1���>�O�0fOʾd�jy
kٛD����ͦ1�ߴ�?q��$�?�}�'��(1n���ڒOU)Ss���Z�[���$�^��Y���ժ/mkQFK�(��I�HOt���'��Ɂ]��Z��JV���p��T�ڰyFjI)ablA�	۟P�	ߟ�R�����n>q*�@�~�B���'�1'�}2�.c����%N�h1#�%)���P���/�����Xj���*�/E-3CR�CX�%4D��囍`^��d�O��d�O�˓�?)��ET(f!�u)E�Ԧn%t�2�mր�y�,B C
�\)�	��jST$O,��'�����d�+U�P�o�џ��ɎS�ؒ�������dڌL%X@����z�A����	�|�⨎�r����f�|I�x ޴:�8��j��_��$ �gZ�\��P��	:yv��z��ɇy]���gC�A��"� ,� �b�̳ZO�\��3O�`�c�'��Q�xѴ�ǡ-���FW�#�te�#~���џ��?E��G�
&8�SH٢ ���[5!���x"�jӜ�Η��ӄ�C��c�;O�=E�d���ƐI��C�����4k��yª֒Q6��F@J$���@M,�y�.W0%�%PF.�=N�2�"�e��y�L�D���i��r������y�ǐ9>�N� *��d�bdU͏�y�CW![W�Y�Jt����e�R��y��>0���Bh��YO�9�-S��yb����TEig].X��8����yb�2���SN��9��I3�y��P�B�	�#?�������yBfL�6c�ѱ �R,��ytH���y�ο�̑��$E$N7�����ý�y�,��u�ҥQ#�S!6�f�X����y®KC�����I�:;=�p"E"�yAg�DZqBD_>���Q�C-�y���5jж���nW�x-��JŬ�y�D �����˛P�*�I�lٯ�yB�ݫc�-+f��6ux�12�͹�y���jx�I"�0~(z/W�y��E:>`�9�V���gK���yB)��D��@��7T�9�6e0D��)�6��(`qL�H����g�8D�<(� ׁ60���ͣl̞��1D������HB�L�(K�aʱg1D��ѤX�vh ����C�z6c.D�8آ	3�Z���A:@X+"S^!��G&]�!�UH%	����"H7?�!���?~U����%��R�X	��)PE!�D�&��Q ,V芝AP�P	X��m$ELJ�@b���De��q��<�� 9?��#��-��Iir�_#{A!����i[#M_"x�ڴ��%6� �#��uR�$�����\`'Ҡ�p<�γeX]�QJ�%NTV�pSaN.��=Y���]%]�@m�+w�����5%l	�Uh��ѓˎx�!RWʆ�摳��'~ �e�g3�P2�N a��9��1�O �q�"�`c�Oʩt�Z�B�' �ð=9��J+�bu��-��0zC,;}�l�!��L�{`0��w�	�3�␓w��@��?�����82��%��8�1xGD�;:N��A�1'��D*��;o	�O
����K"}o�e:�'�']F����x�ኂ�0�	sn�*���Ʌ"R�I���R�4�6�� ˿�"Ԙ雠^N �K����q���@e�$YP���~|X�;o� >�$�SdQ�EEj('�h�'ɠ`���V�n�|���4n�z�f<T|��V)�zK�IQU�։W�6��ۓ$���%p�f�aG$ݯ��($�xB�I��j�S�@���h�F�[%�ܬ�pp�Ƃ�3bH���.|O,�:'�T�^~��Y!��@��|���K��я2H�`B`�۵�J�`���O��Y8�� ��C\� x��LZ1z��_�)�ƣ@�<آ�9��$˸F����L	^�2��e�	'R�!� ��93�ߠ�J�`�Ǖ�-����'�7+�,���+"�\�ۦE��*���{��ޢ�Z� �{��-h�a�s		�k��d3zpH�	�y�Zcl8���3m�`���o��DsB�<�~R� 1��	"�	�Z?�x��o�<4U�w�ڹ`2�1��K?\O�p���z������,n�]0��^�<��푺+A����'W�P����<��Š|��/�$� (�P�Ąa*bh�F�#�p>�%�3K���o
�q��̱3�TL�'�D�Rh�H�"�%[���>����O厜��j�q��� �F�EU��r	�$R���$I@~5�я�D^�5�LaΓc�0HԎO-}��TG��"��n�	]�%�SN�nʭ�a-�Dc����Q |u�%���
ZV2�H0n�Y��x#�̂�b���׮�0���Z��8�:p5��X���N,�(�ʬ>e��C�C�����<" TA"�']:X�	��T�.dr�!H��4������z�%߮W �����7��]C����\����u�j�8�x��0
(�u-Ό���+h�S�vHp�cP��EV�局��:v���ȓD4�d�c_� �aS�π To�HJ�<]~��ECP�I�EZ��S�t,�izg�M��u��olU ������ eoڏQD�Z��T�Fmv����^k��T��X'�ӝVVʓt$�'S~� v��l�rM0fʜ<;�x�@��Ĭ��Ĉ	3r�7mE�f���R�$9&���ē�8�-�#�&Q�҇K9&b�J$��kyB�:��X�dƌU��{$�i5�Պ�EZ�)�`R�b܂7��ɓR+I�hڤʓ��OmkZ���U#3 x�Ec�������V0&�����T(�8Y)�A&#H�qg`=|�X�A��۹"�ax��C[��1��<ɠL�q{��A��<& t��鑑��O���o�D��0��0��R��ij��Q �1�P'+D9TX��A�֪��D��PeP`��|Bui�k�4�~����G�~eP��F�x�t,���'�|E�SE��T��sDע)�~�����ʝ�4T�P��<D��Q�ƅ�"g��o��*���č*S��|�3!�IO�.���fV�D���Xc��<  ��@�B/�?I �?�Ɍ�?a��
Kyri��s���������y��P�I!����"� Mb��4�ޙT4��!�M�*r��;��D�1��D�H>9��';�E�,O�ɻ��O哮je���M�hO��æ��&ԜGz��L�r���I�.E�g��`Q�F�/�?�Ӏr�T�xE�MEC�0�tM�Ih*A�<��l�U?�O�)N�擶UP6�tփc���8���-y�47�w��xtDX�\��!ǋ-+�g��M��U�e��>e>L9���#-B��'F��Q��ck�=�O�ɗ��'{`��ƼO@�(�/;��X��~K`�T���'4�$OL��I� ���-Zh�'K7Fd(�Cr��H~bG�.�QD|B�)N��H��B,w��Y�!È5k���5�Z� ;�Of��$�n�O�Y6M�Q��B�L#bѰ���t�F�Q$�s�D���6��	���5�*�S��	LJ�xծ��X�?!-���h�$f�d�hSӟ�����ĺBfP���
��f����P�0��U�P�4��d��D���`tjMw JU*�>�d�6}��d�"mH�]$-�"dI�6qr&_�jRbH�l�ho���4,�Nܓ�FjwL�ip% ��6jF��d��6g���OQ DS@�`��$�m�t� {0e�����6��\D�����CY�(k���!�@��do�!��'��̉�e��1W\Zy"��{�1OJXS��0�I)+JT�I:#쐤�G�:�`=z�F�)�p5��c��¥O��K��1УL�P߂�r�r=��^����'�`���'��I�P����'+U�����J!V�l��B�m�8$�=	%��.��Y���^��p�u�P�R��������*�s���O����B<�В���N���{rg��g��t�� W+2�CF��V�{��[�!� r�*�=�p<��'�P� @.�}ӆ���T��~���4R���{�oʲp�����Gbi��XB�A��h��ɵ��H��$�a����/-L|4�_0ǲ���ɷV��	��'��#Y�IC�V8�Z����x����0�ƋW�|�=� �R��%�)�~�<M���_a1i��gV��Zdɗ8`xl%�1�C��'�l$�5�S�(�qxbM��|��y�F��x���Qh/~(�q ֧�?�c�\A�V��B<�`|H�N�צ�ɧ �(�1O���g�J>O�I���1+*�G���c�Z;~��H���k�az��Լi@yb7K�5`�|�G"���H̙��ǟ��f��0=�f
�"%���Hشatd�����^x�����¾*&@,�wN������P�U�����	V��p*񉖊�����[�3h�5���<�	�Q�
���%L,�q�t��!�-:�CPb�"b#l�$��t0��oP�U�G�Z�|�T�<�C�J�<��UA��^'�����JU̓vFXRe�B��(���Ɔ�!����f,�����x�l��	�6�F�>Ab�
xz��k �R6�����d��Ⴃ/�F�*�b7�Kh���x'�
�Ъ"h�ѷ,��g10�s��'���Y�0��h�!�ȥ/mʕ�f�E,�Q���'��ӒK�.0(z�d�5z�	Y@��/
�"=Qo8T=L��
�6�-"��f}r�
e{������}��հ)W�R�ϝ��m�
��� gxe�0�,\(��3� �\����XD�%n��;��]��i1\��	ۢh6�lQs��+�ݻ���O�XB� C��%*g"��'�Bf�G�dN�2��xV�_&��3�I�L��\q�d��?<��ce��z�v��`d�5�p<9��Y�Qf�ؙ'b�asQi�0�<��֊�C\lc NW����8��O���j�;E,��)�l;`D00@
c��H��<��`�'HჁl�3�\8ǆ�]Qd���  �HO �A2��Y�.�a�h�nu�EX�̈WVx:�� �A7t���*���l�'�v�k���)|�u�Ǩ��v��]wq��xT�Ҩ�W@�4]��+�N:U��^樨SH����)�F�D~򆘬r��03K�|�pr"���M��ߠ�&a+���<�Dx�v�Ѻ�� �y�'�4d�C�$6��$2@�]�q�j��7@S&~t8��]��'�����F�:�P�0�-��ۖN�- hժ�(G:"?���ϖ,��.J�A��QRKL�?�~�;�P�
��'2� ���l��A�C�hV�N:<�����	����"�U�'Ѯ��=^���zr͔c�5K�ZAQ����/�>E
���!O��P�>�q�Ás�<�*MY�B���!W�dF�"�m�`�Z&�� 5�]�N�td�ɆJF�4b��H!������O:�ѕ�"3�|=�1�Ӥ/�f����E?AtP`�r�ǳZ�,l��c)|�^�@6hW�i�7�O"�4k՗?�UZƊ�qj�L�U�I���X��0�3F��)5��ʾ�@Y1����u(�G�
9)��;|!���ڞ\���o 
�x��G��a��x��'~V �D��;<�0�ĝ�� v�æ���c���p�׉Α��h����>H�S� O��j0lP��	�=�I!.vr�����e�"��U*�x�f/�>}��S�!��a�H%ʕe�'�@ d	Κ:���0i�s��E��'��Փ!Lȧ	���@'Z.5��f�	$ ��mQ3K�a9�ə�&n���y���6u;�HRˍ��0>����&`\{�N+ܺ�_X��"���<it&�8u��;t38�Q؊3�^�r%d�:[ppH���x�����I̐5B�ՠ���<�Fe���K!t|�OF6-K�f�n�Y�B �:����¨L�2u+�柯a넁��g��M�:��u-�9�xBL�q�'��-���E�5�$9#�"Ȃ(��!�bIc`�N=1�F-�edWL��+�$&vl��aĲ���s��a}bHad�^��'q��������@5#iQeY�'����X+�"���A��	���$�����f�|R��J2��iz�c�*	F `�!�FM؞���G�%H�E�_$M��WV9g+l�S`���O�������lJ9Zc���0��lᡬŸ, �dNCEzi������ɷ�M�	� $�e*ڢG
(=A$-�B��2I�صC�"HP�3e�E�!��ET�M�b	�;v�f��cY��X�1�J��0=�$A�@��̚S��0xܰ1��*<��Y�b��<���r���8Cp>���˔��M�c�A.4�a֗������^i�I�A�W	�:���9q�R�S2���<9u�B������:����Xx�C�2��ԺIf� ��@�}�0U0�%[�,̬�blN;Bz
��$���vI����uڞ}Ƀ`I,Sڒ�;5e��K�
PY��ɷ|��OVhx�)�����4tD�0��PSK>��Q(�	S�Zi�ȓ�hɃ2h=8*`��#�ާ���Dx���&1c�	x�`��'�·T>��兆q���D���\Z �ǃm�鉣�.,���Ѧv��Q���X"��e&�f3�y�f ���̓O�x�b(��?
�H�a(��r`h2�$P�d����i� 3!���o�yZ1O���g�39��KRbA�{2�DZ2QQ�KS�]�b5�ɫ�mB�\S�$m��t%��(Rˏ��p=a0,�yB1��!�+Lh���a�3FC)�s(��2���nOx�(9�酊^��ik���8`��&@�i�<ɗe��'�n4��o�V��P)֩�p<��S�-�Xd�wjP�'�ef앚S}�IĕN�.(QVď�=a|rI��f�͛�B݉MT5)�M�_�$�za�ʪ]����@T�F����JB�W����cJ�O�T4+�	]�!�O��#��!*\�)�F����	7E��X��d�7D�T��	CI>q�Ϗ�;Dv��#��
s{�i�3����B`K��|2��r3/�4��
ۓ`k� �W�O�.b%�%Q^)h�28=��(FA�T⑊V� ��S�_�P-@'�x�I2���% t!%Z��P�W��U�ʛq�<ac�۴!|@!��<R����v��Li��F�����:gn� �ʖ�lac�|�R�����cd�Q���4�T� ��=��[mX��;��P�^�<ȱ�T	b�����T{�8�pQhʂM�X�bR M/;5P��,W�-ڴ�D)"����$��1h�J0�V����R5b�������J9c����BŨe��YsʟR�v	�-���i����'o�@�zfc'$��+��צ!Q�qb�W��eűD�!�DΣ���i��D:�|�����!�$��D"�2�6*8����H�w�!�dƯE�4Q$㏼l��0*�>B!�I�`�0��M�8�j�CvI #{I!�I�$��4;�X;�Z��WG�&�!�� 4hp��0w���G�"`��f"O^pr!&� E��UW'�`�X�"Ob�����{7���oO51pbı�"O���GJ�@�B����8'n���"O����:�j�P�K�,-Y��F"O�q,lF�[cB��;� ��b/>%!�dݫ<�x�j��кeh�S.�D�!�$G~'8�bvBϪhY��Q�|6!�$��.����%쉃EIR�	fm� >4!�T4~�V��	C�r<fJ{�!�D�1+�6ả+�"�.1	Zɂ"Ot1a�31��8�Iԉ.���"O���(�20f$
G�_<!��%��"O�dB�!ʜ���FiO�Vh@��"O��4��;&� ţ3�T-�"O�%�vG]�x^���gP;	l�@K`"OĈ����<����N�eV��Y�"OVa	U�F$S\�`%&�$�p��"O���+G�3�v�(���YÔ s�"Od����3$hm{�왳~�ʨ��"O����.�.v��R�\�~`�5"O�Yv�L7mt��˳�E95v:-�P"O�� 1n��w�h�Ϛr�̤@�"O\�3GN*Ո��C#o��=��"O�5���i�ȹ��OG�TnƜ�c"O�(0������4�G5cO��"O �&�d��Dx��j0�Y��"O\i���6�Vt���1Ǧ�B"O�0�w�Z!O��(�B�՝�z�!�"O�����8=���F����@p"O⴫֣�:N`V�����l�,L"O���l��d>@��1q�D�4"O��C����t���i�a .�ܑ�A"O��86�܏-�l�2�ڟx�V���"O��c��VÔ��-�.o@��"O��r2k��<�p�B̚�hT���Q"O@:ƫޜ|,�'�\�1ۜ��"O��rT�T�b5�P2g��=1&t�*O�ypV��^���1�,V5P����'�j�Q3�p�fBB��Y�'R��ac�:*��=0����wm��@�'ܬ���P� IȕJѕn�r���'�$�Ѓ�>��>Fq�'ܢ�c��>u���A�2����'�>�p.15�T�iō��%��T��'�6k0��1Oy(qoޠw)���V"OL�"%c��A�X�P'�'1%�\�4"O�`IQ)�*'D��Ä@]1?ji�"O�h*�MB�0�T�F�R'\�0�"O��Hۘ,�v��FG�4�f���6D�d��)h��(��G�F*hBF7D�d3��	j�����C�A4	��4D����3������7$g*�x� 4D��(��  h8�}h d�vy�2D���@N�.D��P���H���ha$D�"���_��ba�F T��7D���V�.rҤ��ɯ�Ā���5D�DX��ޑl3xmYWȇ�FsRrE`>D��R��-�\�y"�6m?
�Y6�:D����C-)<�$�0l�f����D+:D�Tj�4�(��".�
x��S�9O "=!3�B�%���FC·`�����Ȏb�<A	J.:��<���(D��Ժa+w�<i $9-�X�H�آ3Ir��a�t�<� �.�����P�'Y�k�݈�"O���5�USl�����2���iB"O8���eƑ3��3�i�;eY����"O�U���4w^�AFɝ28�l��B"OZ����t��u-�~���u�D0\O�dp�
�G�h�aO_=����"O��0@Бƈh��NQ�h�q�"Oօ9@+ѓ��5����8�V"O��FV���YՋ�8w&���"Ox�a+�M-T���N�0��"OI�T	W�><�i�D��;�8q6"O����s6�� ���T�K "O��zq)��T؆옟_��y���x���I�	T�$��C�G���	�k�+�!�D��v���@�Y6^�6$rG�O�!�d��!�VT����%f�|R!�J'W�!�$.�5�e�<pyzá��[�!�I�=uFq�p�� QF�
���L�!�D'J��a C%	D呵o� �!��ҴU�cA��>�)P �3 !�$A(�~]�R���10k]0K���M����͢����T �+Z(�jh�v"O�9���M�o�@���Jŵ���H�!��J�9�dH�,F4
�� ��G-�!��SvN|R���*:3`��r��<�!��?W��Աa��nIJ ��*�!��ϭl��T�H�)9A�a��L´3�!�.[�� �6�� 5���m^�G�!�DH�z�@�B��z_V�!���S�!���C�ؤ#�һC2)��&ע#�!��%�� �D�S�+�Ď>Pi!�$ۅq.`Is`T�O��Ȼ���;l�!�ԋ�0���
44��{���^�!�V�P���2bZ�~��g�N��!�� 	f\4a��%d��1PA�	k^!�K)=OF�Ҵ��d�ޡ�p.�}�!�$C^cV%�t�Ҁ:���ˢK�^�!�!�R틧f��4����λog!�$�6��(B�jXx���)0r!�0L�FHz�� �28a�[�^�!����M�M��S�.�|�!�@H-N���(h,QmF�x�!�S�H�측���<P������t�!���f�i��d�: C$aC�Hn!�d�/{P��CoZU�,X 2E@*j!�Y9;�85�e�r�m�&�ˑM!�$�fkh�RF'��e��u$I3!�ۑªa��
D�7��2��?/!��Ӥ
��4��UY�d�e��?y!�ĝ_p]"a��S�u���E�aaR�OP+�偙M�,1�%J�V���"O��Ga��<�R�hgH�
��Tx��'b�ɨ0k��q��"[��TJź)�NB䉟fX��p�!��;%����cA��B�T���%�;2�x6*-e�C�I*fm����a�\pXP�:<�h#<!�0���*�)� )s.	𷋇�^�ȓ#�����RB�-R;*� C剹�Hͫ�+�.:���!o
8LC�ɏ:��(b )DT��� �e�A\B䉈T�<0�éúв�;1��]g*B䉔���seE�;wv�pvg�%u{�C�I�G��0����2)<ᢀ��F���Ɠ8h�K�!2O$�r���%h���S�? ( �N/t�� 	E1��Ai�"On�ʢ�ƪ ^�¢g%�z�{"O�L��f�MJ�ş���)"ORqa��,8�`�]7�h�8 "O��qD�XnD��%d�/���"O�� ��-Ǯ�A��׬7�T���"Or��0��;�Z�k�0���B3"Oډҳ��6U! �����UoJ��"OX<�T�V F���G�9
�A"O ��W(�9y!��*s���_ΔAI"Ob����97�<�����BU� �"OnĲ�jB�zg�0�D��(F8D4�"O�8[�E��~_�� ��G!z"�8a0"O�q�g��o0)D�X�x�<��"OPd�����HK��^;?c>Ps""O���U	V�"ӈ����sG,Rs"O�b�G:8���̓$D:���"O2Y+S��	�֠��M�)�ؑ�"OLԀwA������?�<(F"O�� ��:����?D%� "OXP* gރ*T�e	�kV��"OzY;����#�4��A�P�pB }��"O���] _��H!� �F#\��W"OT���W�D(��*�e���"O�!�Q��/7�p���J�c	v�:�"O2��t%Ó�Μq�IяY�� k�"OpQ�m� '�~���/��Ls"O8;�F�`d��퐅��`��'�Q���]!6H��qd��*�:ea��#D������,L*��a	
�,���"D�0�$���-�f�3���%�"G?LO<㟴W��a�X�Ʉ�S!u��b�/D�(��ƞX���Q!P���Y�+D����Uv���&Xsu��s�+D����n�yl�(r�i�3DP����.��<�OX� �ٟ(�V	y5j��Qj����"O��08<\��Q���dD����"Op�ٕi�dy�]ɓ�ֹ#V(8H�"OB=� ��p���j��<[pX� �X8�Ę�+U�d�!���*��X�3D��.2��Ag�C(�
@ ,z��C�I8V5�x�m�3����C�	�"[�tR�C()�����L����B��>}��R���+��]�G�ϲR	�C��#�q�EB�^9�]�D���SՠC�=kLR5��i�()����M�Y��C�	�a�-B��,+td	p��?C�	=X7l����)�J y
ݓd�:B�Ia���(�A@gM\ᛣ坨/м�=��'v�ΉQ�R3@�22,�5U<N��ȓ���ɵLƅ6���gV�}h���N���
��E ��]RU �$2�u�ȓ��bÄ��`.��ʚ�lm�l�����v �s��|6����K�f���hO���Iϲ~��	0�Y$N����sa<^!�D�T�z�C�J�`-VA��a�!�$�57C@��q����ؙ�@�>�!���>ʔ�cխ]�k֜���h�W�!�dH�3eS�#�aʩ���:S~!�ѺEL���*@5�P�B*�)s!��=�h0�����i� \��	R:M�!�DכD��Z�, xi� ê�,�!���l�J����~Jx���C ED!�Dݑ2���{vA�)I�L��B��@!�� $x��(!�@�R���s qp"O��0�ePbLQ3I7'����%"O�!!2R�`����1th�1"O���b��
��w�Ь`J��a"O\����];N5ȔL7h���"O�)jc��x��0��
�\��iC"Op�F��L��X��e��(GV�s�*OT���M.O�V�0�O��dט؈�'	��K����['4��E��:R��U��'��(�CZ�i��Yf��Dvz���'%��*%�ج~N8� .U�$d�'ZZ�f�%��se�D��� ��'�� ��d@�tB��b$	Ʈ�i�ʓxpL��P�!�L6s�����i�<	��O�"����9oj�QH�h�<�A���J@%��4R����VK�<���_*�:���gD��
�Xg�\�<Y�kk|�q���V�L]ȅjQ}�<�c�ƴkjZ����H�.i���x�<���~h!cQ��a�`)�eRt�<���B�ɀM"�	8d�M��"�l�<!�oѻ%f��H/&uaƀj�<��ㅗd�~�C. C��	���^P�<10��7_�4�bi����T �J�<�Ek� �x�v.@�)!J}��I�<aw(Y�H+9��`C.@0�8:D!�~�<A��ٸ>,sB瞪U��4����w�<Q�#ܩ0�N$�v,�6�4Tv��Z�<�e��[Ŵ��Vf�>Rp��'�W�<)� 7�r]�ċ�~���ñ
P�<Qp��-<��9�Pn-�xk$�N�<��^�;}fT�EOт  Ph��h�s�<I�%�/�lс2I�>41يBg�p�<9�[�VEv����z��]*���l�<�V��/��01&� P��ԁ�|�<�#�I��0 .��m���-�Vl�ȓ�ܜ@feÂI��,�Sc��i2=�ȓ"9���*܍6���$�[LnM���Ā�`J	f��Ha�i��V�ȓ��9��W�9����L�e`0�� ʉ��䛮�j� ��� I�Ҍ�ȓZY�ЀOP+r�X@5�%m���V�,�#O,D��;�#�è��ȓ#  %K�� I"�T	�n�̜��ȓ��0�LZ�K��Xp!B�4�2�����e�y$��1DX�7UH��'�U�<a�L2QvL�v �v9�H�k�<�A"�&B���!jˎt������S�<! a"L�x���J	��`�ӏ�L�<)5�^�>�%�Q��gZ�k��C�<A��I7��P��=+HkŁt�<��vx-�fk��Y�Vqp�z�<�0H8PӖTEf͢uo���C�Ls�<�,�<Xl��ဴ瀠��I�<�5� Ɍ�QJ�n�Ș�2L�k�<�v��r!0d@��I���/TJ�ȓm(u�i��)*���ǰ.1"(��3����GO�Lo@�iê}�f���Rf���q��1c����D��U�¼�ȓ��a�eO���0�bh��f*��ȓ>�eR�����ҥ�x�&�1�'��9TK�p�B:u���s�^h��'Q����<���Ꚙs%2�*�'�V�I�b݇%����w�_�>�J����� p��&-˷`H^�bfiY�03"Oxa���>)rH��"?����s"O8p	֯�l/�t����/a}���"O(�b�J��Z�m-SnP��6"O�ي�!6!L�����T.i��c�"O~y��BJ�
 {���"O~Q"m9�t��
�.
v�8A�"Oz,�@e�%�z�{bg�$`�y�T"O���"I�3<�$��#��)<�a"OT}�ѧ�~��h4M�=Ld�0�"O�Ҫθs�fx�R��8. ���"Oؽ�PN�-j����	�N,Y��"O�9[�]<��ձ��I���!�"Oj���ϩ)�<`ai�4*�b))D"O���g�0�2Q��_���z�"O�9��� �/�~���G���\3V"O���f�5��WM`#��V"ON�R�	K^�	:,ڮQ���"O�D��T㆝RҪ.}�XIp"O�ej�9v����3g��G���"O����\�J
�I��ƳG���W"O ���7�,=�q�� R��Mچ"OԸ�	Z�V��&,�1�\U��"O"�RjF�d#����Ѷ/�b�!`"O����I&��Y���Y���`R"O^��Q��4p ��p%�&!���T"O�=��g픤J�@ȑt缑["OD��	_�{!�T���#�'��e"�YuB�R!/^��@Ahb"O��P�LW�'4hI�䑵��+s"O�Y���0>��!z���Y�b�Rf"O�0�$���0��H�_:g�59#"On����1�b\�V፨�h��"O�De�5�6��ρ"6��̩�"O��J���,-L@��/�>O��QB�"OtuH�*�.WN\Y"(�(m쵨"O,�X�H^	bF�1p�5	��e8�"OVi D�e�(ʃ�
�p�$��e"O��
K�,���(�[��&Y��"O`��pI�6�^]�P��&�pP��"O�Q
0(��@&"���'�?Ihd@��"O6E��oI�]����OI�����D"O�=�럋l��ErT�!�6�Ӵ"O�IB��SK��u�M�M2�iг"OP�H�������Cn[�y0�X �"O���mQ���8mD	j(9K�"O2�3tO�=,vM�C!�/y \,b�"O�i��k��d@3�6m�]R�"O�!!&`�cm:���KK�``�P�#"O0��$c7��E$���"O�P!����*"����ʆ�IU*�[�"O����̂��99%j֩M���"O>��Q�\�Ia|y�(Y�5-��k�"Orx���ǌQ�" ���2��"Ov��c����X{�	C�~IJ�"O.!�wo�6=BE�h�]?��8v"O� �.}�8�s��V}*��7"O$�x�!('�۴���dH�eB�"O�i�6j�	V����ˌ�(9�pA"O<��$ғ^�duؖ
�yV@ph�"O����%�qT��hQ�*:ȭ�F"O�dR"%���4S�eʜ-����"O�T�Db_ ��q��eʒL>(���"O�͡"n�N$�T�ʛ4U��"O� ƨ@7�іf{�Ya�Z�$ek�"O��`7#��
�8�hgE������"O��W��bژqԃ�!;�,H�"OU�p�ֆ_G~p	��)�ܡBT"O`�8W,5)�	 ���
���"O���7�Y�{����,^�An4���"O���m�29K�F�?�N�"�"O��PG��u͹�*Z	0�,�"O,�xE(#m�@��'3E�Qb�"O���.NcM8�2%a]2~���P"O����Tk��g/P�u�jC�"O%I��γ3x� ���L��"O,�,)�§G
.lLRUR �6�ybk�r��0X��R�mb^�C��yr�M����:�&�{MT�Cr�/�yB��J�& ���9<��q���H��y�F�>9R5�V�3Z��ߋ�y�� 䲔S%iɾ&�V��`���y�fM_,j����P�8�KEd��y��I�0�aP� "g�� e�?�yb���|Ę��E�	�f!�QRQ�[�y¬]�0R0i�Ysx)���yR'\/Pt����Ĵ��T˓�޻�y2�c`hܳrK�]
��CI���y��ÌiϤp(6�FNxq����ybB�8U$u�B�ԦLv�uY2Aʓ�y��
?{�8	��*B�PѨ��V0�yR,��[�N��V͌�ܖ5��ʚ*�y���1�ԸmݼbRT!���y�i2��RVo�-��`�K��y��WJ��ؐ0�� T�J`hN&�y���v�f!�C7Oa��(g�Ǎ�y�,�x@�5{���L�~�(�"�y�oܙe��M��^A�Q,!/��rp��S&T� ����"Vҕ��,_�x���@���`�
�6l�D��vfR��*�i�`h!��)p䉇�G��E�0G�F�����DJ����@$�]�E!�a,� ��FT�`�����rq|�wL�$XR�ܲ���5u9���TE�`�ۂ=�jl*��DL%�ȓ^$H� R#�ҭ:�
�&�P�ȓ-������ b�X�n�<��܇�x���G��"�J]2���5n�d�ȓ��#��'_g�݉��B�K�8�ȓT��%�fmPN�T �CQ�ц�l�jX�$�g�D ��X;nM����n�6�i��
4��0t��4KgXx�ȓe�
Qx�Ź:F�Ȅ�M4f�C�I�9r
��2�?4|�s�'{"�B�	�<���:��#t�8Q��S'{�B�I��H�  oy{&�h�=i*�B�I�$���J���a8��t	�	w[�B�
'��Y"׆4
��0=~�B��.c���'S���ȠЦT/y@�B�	�\�h�z��;;��E�
�}وB��2c���'
]�`�<�"�m��RxB�v�:�C���$ЙJ���jB�ɅN���J۰;�����D��C��C�L<1��!Q� r�dkR�8MxC��=Tb�*�c��h�k�>"L�B�I _�)�sĐ�%N�рNW�s�B�	Bb���3� �
�GćKu;�"O,��u�*Z�I@ze�"O� .�)����j��#�_:���"O��Z�(�]|K96�1i"OP��#ɑ�Z7N���"A�a,A "O�@����X a�R�:@��"O�k��� \0Sި90\�XP"O��S���SD��ԁ�/"V��$"O�QTi_�OBI���9�<PC�'�1O�� '�-w�� �IO.9�\�"O��Q"��LM�u�W"��~��8�2"OȌY��T�Z|
��`�v�a�"O�	J�X�J�,�����zh��"O��`��*G�pFc�3o>�2B"O،�6`�*� (������8�"O�xPF)�:f�*R�IH�mG*�5"O*~x���Č����Y�"3h�!�:f�T[��93�2�`�ʩ�!�$�J�#UQ%|��& ۊ �!򤆒=JTP4��#C������!�$W
u�Lx�R愔G���#��X*an!�DD�0���#7��E�R�_�P!�Ē����%��2Q:�-*Պ�/�!��M%=�Pq���G6b���#�(�!���d�����e"6��"��!��؜x.Y���7^�e�d�A$%�!�$ސ>�86C�]Y|1*s"�/XB�I�(]�9���N6��&�s�`C�	��l�q-�B�De���9a\C�	.(���ŕ�7E�	 V)�/z�6C�I]���{�����d���.�V]C�	H���
��,��I#�a��m` C�I�&��J�"W�q���PH��q��B�I�c(H�A�]?`�`SC��LI�B��	Gy�ih抎9;��l�H��[��B�ɮm�4<k�P(���Yg�Q2�*C���U+�&`&tt��AմK�C��U��!{T$H�q��7���	�C�ɊQ�2́�cG�l"c�P�F�C�Ie+Ζ�&1R��'쇖����s"O�B4�Wp ��Q����"ODq FC�s��t�Piӓy����"O�a���I/~x���� }0<*�"O���� C�v
��� ػDo���"O�!�@h�0Y���J��Ś=_Bey�"O\UBAl_�#�� ��<c^�D"O*��!l��4 �����Aؓ%"O�HK&�&�hQ ���e6 a��"OؐR���*?��q�6M��t1� 1"O���`Y)��b�ƭ!()�a"O�]���6��\�@A�|,r�{�"O��I!n=�U
�`ܨ-�\��"O T�7�Č��&��(6F��"Ot�J�&ojX)�3ˁJ0� �"Od�WE �1��
��.�q�"O@�s"S��>�KӡY岘��"O��k�k:���a� }>} �"O�)���K���	���a�ƹ�2"OP���DZ�|� X�"#)
xMR�"O�P���	tn�� �K?����"OP����'x'�9��c��S��Щ"OP�9@T�w����[1z��K�"O�E"��
���(f�\1'���d"Oҡ�"i�!��bs�N�3y0l
�"O���6�J9�Js͒4x�0̊�"O��)��e����˖%"���"O� �B��^Mj0��-"F؈�"O����OrC(��ә^�J!Ӣ"O �0s�ʯg�*4#�㋴	 d`V"O�չR�[<�� ��$x4�"O�ɚ��
4;�$�S�]������"On�J�I7m�:%�׮�=�x�i4"Odp;B�S,,�SH���"O�AJ��S���Rӳf��c"O&�2S	T5���5Cʟ�6iR�"Ot��2��9+�V͈6�ǚ���
�"O��p��H��%�a �� w�09"O��#4�A�V��&Ā\���#"O���V�/l 
`�,� d���R�"O��F��sp}���A"�aF"O���FY7;�X�{���8E�
ubu"O~��P��<Atڲ��%`[6XJe"O�튂O�J}n����t��t{R"O:8z����O����q��w��	T"O�A�j�D� ���Q--\EH�"Oz�g,[��vP�G�![�͂�"O�9����v@,TCF�&��,�"O�$X��Fm8�6��n��,�R"O �y�q��q���4X�&=��"O�Hcs�,@@򔲷kL0h�=�w"OP�8��.iPݑ3�*u�"Mj�"O"�:�fW?W�b�k*����Թ�"O������m��h��Z;>�!2"O^)��	�rnX�s�hټ�z���"O�0��ʹXʙ��'�<tQ�"O\U2��ҞGl��g��!��yQe"OD	zG*�28�Qڔ-�j�����"O�Y���L�1rL�=+ڹ���1D�@:P�º Ȱ7FY�*��U�'�0D����	+�䒓 ˱ۜ9d�+D�0�wˈ�He�iȗE�z�va�rM)D�����+g(�4�FBԅ/�\�c7�(D�D@�&�
p���3��+S^�qSf�'D��gJ �Y �m[�IqI4@2D� Z3�C��eQ�#T�`�Ը"�/D���0��:ִ��c�Htv��#�3D���DB���i�f��>rCh�#`�4D���2��&f�6 P��K�>B@�u�>D��SR�ٚZ�<��*�	����n�<I�c�C����	�P���8֎`�<�ըB�#m����^��%��c�<Q�\�RFnX���ÐtVv5���^�<�t��5�U�-�&0N=�У�Y�<�K@6j�����Ѝ?8��BB�|�<�.�"K�;� s���d s�<��c�	�]T��l\��C�<Qr#ՎS�*����u��P�T x�<��n]Du Ԩ�FU�U����n�<�r�U�ڥ E"Ͼ��k�b�<94�)-�pA�F��BЮ�z�<ɗ��/,V8	0�X�w���H���r�<�e�ԁn����L�&>�h�dN�q�<S��U���� <B�ȥ"�p�<A�D^	��<ɱ*�
<�,4 C��B�<�'��s� h�
�wb(D���I�<�!W ]f�ED�ϖG�B�FςF�<��䌳���H�D�`�4�U,�Y�<���W!l�J��%�����%dC|�<���Vlr��/�>�8�z��0T��asC�mnQ�VA��\f<w�)D�� 0���I�;Nn�
�D+e���x�"O���Ue۝eb�Yb䬇��qZ`"O�h���'o��m)f)Û����"OʀaW.K�`�T�vO$Y�"OB0�De]4b�1#-Nw�mp"O4h:D�a���Q��F�4m~h�!"O A���_͘h�B�XW�D�5"O�}AS�� �d�h%nG."Æ"O���dE�*BKEG����"O��5�B-;P�������t��w"O�&��j耕��cͷh��Y�4�'a��^����PI�����!�$ܦ2�^D��aߜ J12W��!e!�ě{��� ��?K��<`�)D#^!�DZ�-�x0+�h<�L����"A!��#p��4X�M�M���4W!�9G�;W`��	����'���/!�DA??� =0�Q�X��"�7	!�$�R�̭:4n��$�`�A�Y6[�!��p��ikF,C9�6�x�l��g�!�$w	����)*j�� �T�}�!�W�>D�� fo� G����5U�	�!��}�z�J�����C�e�0O�!�D
v���SG(:�3�v�!�$½�����C��~#��!�a�q�!�d�=��,��oڷFUց���!��>]����GaӶ-�L��D<JU!��$N��ɱ��E�����A�!#T!�$܄
묍HÊ�nZ��ce��Ag!�:DB�<xe�E�^�B���'�!���/P�2���(��������>�!�_Y�J�� #H�%��FA�v�!�x��w �^�ti�ӆq!�� PZ������g$����C�Zh!�d[ {W�]�O��@ �^)NX!�DE^��Ug٨$�`D",33!����La3���8#�f�4��9#!�%tt8Ҡ��6Ϭ\���	�!�$>�BP"��٧uͰ%��L�v�!��+��|�e�J.c�lp&e֌2�!�C66�2&HQ�e�B�RMN*!��N1>7|!3A�ۅ�H� E��'l�!�ޝ]�`�R��%��t�t�ŁF!��:��d�Ųwk�`���O7L�!��%M��K�m��{X�h@pg��PyB$P6i��٪ �.$��s�±�y�*ȗp�@����.}��S���y2�^��\�0�H�<Ĭ�����y"��07 �R�	��u$Q��
��y�'�6L�e8׏���P�h%!¦�ye
�g	� �ҙIcv��DDI�y2��8KO��B-��+�Q ���y�연Cv�50��C�)�2�� gR�y��ȵ �"��3��"4,P����yB�;FP�YÔl�0��,;`��3�y��H��-�e&�(w��( ���yBĔ�^�MILDxN �g`N�yR�N�'��4�)0Bnq��*��yR�.� �)�b 69���PB�.�yb� �h<)����U�9�@���y��ȡ����D��n!�����y���iu8HR�ò`?�Y�@R3�yr��00a1ǯ�Z
�������y�e�m���I!"�}#�Z���y
� ��Fc��:���4L�Gc�Aؐ"O`��4�Ѭ%g�$�
X 2�UBR"O6\��j��q�X!d.�9�"O��Ȣi��Sz��1F)Յ }�"O���:,�(]�g�XeR�y��"Oj�pQ�D-#V�(Gř6,����"O2"D�T;$�Ex�B�_)Qc3"O���S��(_'�|���T$C���g"OZ���,k�¸���A0S�2}�B"O�T�׭��m%�9�s&�o�~]#�"O�8���#nye땢�!�HdX3"Oqst��>vT��WBF�����"O���
�z�s�&P7�����"O���O�O�Y��_�B��"O���R�T�TE@ؑ��(Nhi�"Oz���V�+#�R�
�� ,��y��֩ �6챕Ġ6	Hu�!���y�f�2�����`�a��	q���ybO�H.,D�����D��1"@���y�S:BV�QMޓs)��"&ך��<q���	7z��dѻv����a��ax!��� S�Y8�F�8���A�-�'B!�D �R���8��hn:�{PX8&�!�D�6l���!�MO8M	��"@,�2)!�DM�H�,�S�k	/!�:-I�
J- �!��Y�p9:�(��慲�oƲ�!�O'"SL Q�o�9*ф|�.5�!��]�kuH$�բ̏'�>����#g�!�dZ-(N ���%����"�ߖ�!�$�/ٮ,���)�l���D�88!򄇏DS@$Y��� �BHH��>}.!��8��`�.#��l�� �j*!��(.l�S@�10����� 	!�ē�{4�a��%k�@H���*�!���*��8kf�W�O���B���H�!��XJ��I�	ڇh��5AV�1\�!��~�j�$a����W�O�!򄝳9z� Ŭ
�'��XrQ�Z	p�!�$�&n]�|�Q�	�|~ePT��P�!�5Jq*T2���Hؖ��*N12�!�d�}�����BٔD�zs���j!�Đ�J�`��a�,3���ۅ���vS��$ģtD��p�� ��E�cG��y"�F+aRNY�tH�vjH4���y�n[Jv�R���#�� BR䉮�y�l�Y�5�$���3�I��#�y�
ǝ �|��H��3�Ę�yb�]�&��-����J�pH���yb&\�h\�P�?L���5���y�F�m� ��q�].wP�M �mʨ�y�Y 1.H9�`5}��ʑi��y�K\�$�P�����o�4��C�^+�yR/����E��.%jTu�����y�����@K�c�^B�ː���yB�C�^��09��ӻf鈑X����y����G�@�p���R�Li(P���yrd:]8��Q���\9(�N�2�y��!N�� �dE,	�:e"�)δ�yBH �Qx��˧,T��U�щܞ�y"A�<e�Ь�� �`��i)����yR�΄z1 }1����'�X<{˞�y"��M�p�RN�  ���o���yb�qX� r cȿD����+�y����h0��]oNa����y
� �R�"�-�`o�D�̡Q"O�����ߊ5�l�&�O�q�D�I"O�P�ąT[B&�A�,@�;���ȵ"O�aӕe�N���X�%+;~ވ�s"O����*U�4�a5⟭ln ��"O8��oB��X���bW�n���S"OE�G��"hL���_kV�͚0"O�e@��4��8�e.D-�)H�"Onq4�E�2 �m�Ń�36.�cw"O�rb�כk�J�p�X�hTX"O�ԒB��/:�x�����$��"Od�"���:��p��Mӱw����'"O���WF�*w8@H�-��wo���"O���I�?5��<��.I����"O�A����k�"բ��B"Zt�(�"O��{a��+k��%�m�4~72|��"O��F��xX�s��S"X��F"O�	�P�I�
�Ny�
+���"O<�!޽��IrD��3��H "O0	�

I�$X�Ò.3��P�"O$�"��)�=B�DY'o��""O<�X��Va3�	��#�#sh�آE"O�\Yr� $D�*H������Z7!�$���() g�7�YS�D]�<!�ЌT̠�h�F\�L��pI!n�^�!�DR,	�\��!K: f���'�x!�ĉ>�,�#,�Y5r�ゴV7!��1u)A��b�h���`6x,!�B�e,jhA #?J�b�bCOXg!�;&) ��ͣ�8q� �C�u�!�DL6|�J�ѧ�n��T[��"!�"/�f}��\�c�4͋��:�!�d�j$����V�j5���Y�|ǡ��;�2�;nL���'�gIxC䉁1R����D;�8�iBǈ�?�<C��8߰��vet3�4Ц$��.C�I>,�Lyr�Jʷ�椲���)��B�I;bdP ��\P�͡p:PC�I�m8�郑�ag��;Bǉ�b��C�I�:U��	��q�V9MY�C�	�i����.�0�jU��&�=�tC��	'd������@�V��㆓x nC�ɄD �eI� �T�C�nC�I�/�d��F�&fR5�����>C�	�KB��*�GK�,,��t��`�C�I�#�.�1lE�&�.Ъ�%B}UFC�I^�ɣB	��NV�T3�n��E�lC�I! Ѕ0�Z~�\�ƭ�W�$C䉚.-x�dϐ�7e�TٷD˞=�.C䉀
�hHY(� `C�?������3D���qi��]��pcGN+h�+�?D�4	�.�Y��!`À̎h�P��S(D��@��)]���#��=)vf<[�i'D�t��-�y����1g�y>H;��14�<�f�
H,Xy�$�$E�@�ag\�<�@HM8n�8`QT�ޟ*Fx
�B�<��JH���BG��nPB4
�
�r�<��{
��2*����ɹ�'�p�<�r�b\LA���@%P�,q�<�1E&�=)���/Z���s�^x�<a��!B@dM���B6J����	�x�<Qq�UĚ��҄��d8���{�<A��H�xd��K)D�ī�
QC�<�	
�^�R�ۢ-s#UɞE�<� <�(�m�&��ķ!]�-��"Or�p��R�BKX�F"=�8�"O��{T�"�
Q�p�X�61��q�"O2�;A$~����%'�V L�!�"O �B�C�=M�0Y��^�DP��"O�C��\������6J���"O��%G�A�5x!DA�X�^���"Ohm��]N�~ykE�M���""Of-X����pK�O.J����"OFLa�ċ_:����(	H%V"Ol���h�-WN���`F\H8���"Ot�̈?�0�B�;w(|ز�"OX����"㊏u"��"O��J@c�a��y�O�n�z�*"O��a (GDZPU�_�>�j��"O��	EFJ�A2���J>)�'"OV���
m�D��l�
YRd�T"O~����YJ1$MS�7Fݮ`�@"O<����D  �b��*x���$"O�I� j@:gcV!��F.w;���"O|��曺3��L�/ġ[6"O��e�ê9F�f��F3�`ɵ"Oʑ��.ݿhe�9�ł�04a��"O��A�L �<b�����wGބ"v"Of��&J�b�	&�A"e��Ö"OV� WcK� Dj�㏨3Z�S�"O���fN�X ���+þ`��h�"Or����:����i�9#��g"On�'��$c^${��/���2"OV���N��$� ��F���H	�"O��PI��hy5�M!d� �`"O��!&��E��Z[082�"O���
��x�@)X�a��1(�M�"OJը���1��ݳpAڢkr�0:c"OƘ1waœ�l���� zf���"O�U9��3M��;'o?� �"O��EH�k�ơ�͜v�hӲ"O�@�޸��}��ӕ(�ٓ"O*��(ea�\j6oσ)����1"O>�x�͟9�N�@/�$�[�"O�)
�l�w�T�z�퇡z��"O�U�C��3d���	r���"O"��Hع.��=�u�[^�yg"O�9��P��%�YZ�j$"O�B��ۀ_M�)2e,-�:�"O�D$��=9$�����0�"�h "O$D�Tey���C`�MTq� �'"Oš��VD|�ɡ�n�1��mq"O���F5u�~�b���O�D"OL�dM��m5���g��F¢�"O^�Aԩ4=i�b4���l����"O� �Q
<D51'A�e�|"�"O�h��X,ALX���/J,O��Y��"O���#�)3<�X��Ȍ6�zq�"O������dI(c2Έ�
�:��"O�Y�5ǉ6�x�m�I�g"O��5-�q�^�L܅e��86"O$a�Ӡ�2^�$���.ukS"O�ŀA֗+��:�-� }|��3�"Oh��`�'H` t`so�!}�Ԫ�"O
DI�Z�O��@��{pHx�2"O�c3�ߏ(�t�P��(gL���"O�%3�W�?≡"ƙ8DV��e"O��;׭��N����d�]	CD�c�"O� �Ū���%P�f�c%�X;F��a"OD��\�`2Q����l5"O��X��2�H1�5*��Fw��ˆ"O�0�GC������@l���"O�M�V�+8P��T�!  �9#"O��c+�%a��ta7NY�E��"O�{���8����M�D�:�e"O��d�ߦT @�/H4A����"O:�A#��E�:�:��Mz��"O�kv"�/z���&�Ǻ.9��Af"Odt�W���m[�@���Ps�"O"=���E�XHL5�#E�<k	^9Sb"O"�(�(��ʱ�#��x�j�S�"O,�`��H��7�76j�]��8D�,� mh�> �C�S,d�S��6D�@�CN�0P��50���%J�Z�
bo6D�p×�͘M��9�j˺{8��%�>D������9c�e�%	�-�ql'D��QT�H�!w��4���fy���2- D�\)�ڷ:���ʥ �P���L?D�ܨ��UZ,�8�ʃ��@��2B=D��jPΟ0kHY�ŉ��qBy��;D��Xp�֠w"���	O�A9�9D��SЂ�)Q�)���'w�7D�Ă�4SV����V�̄��(D�����8EiN�$��
CԮ�ԇ&D��	3"c��(�)أs��L�+%D��p�҆9�؉C�T��|��"D����!8�N�E���"1|�A��>D��Rf��*O"=ZT����"�>D��	&���6�H��0�"P>��I:D�h�ďW�H�'U!j]d��3�7D�r���$	Z\u`WЀ hJ����3D�x ���z�����+Z�f~��;�7D�pR�nW5b'1�Y|3lձr�(D��$ `� ��M�����%D���C�h������N���!�N1D� ���F � �P��ʎ9Nv-j��0D��V���7�z�
�ɿ`����G�-D�(���ݰ1�8��r(��;Ԇd0b�*D��Z�lI���1M�V�J �:D� a#�E�\���Z�g�%o�.�j�:D�@A�Q<�<������BK��I�~C�	�`8�Y;E�]��<�	��ݤ{�zC� A�t�
���@���Z���RrNC�I	������G��!�7j�@C�I�cF<��%\!x�*X;ש�"�NB�Iw}8��GI�e�*�1u��/j�C�I��^d��C=]F�k#�ZtOrC�ɦk
Б9S��$o�2!H�L�.�PC�	81�n�# d����)"jD6C�ɸS:�3�� ~`�Dp(�v(C�C����EU�t��8S�Q��B�ɒ0�d%: ��L�<Á+��*W�B�I������N�9&θbq�T ��B䉲w4�t	/�Q�aظ.��B�lO$��⌝q�u���֑e��B�I�/�4��JC�196�^��B��/R�Kg��4��y�楝0:,C�6b��(��,S�Tx@�ډOC�	�9��-E��9v  ��gx�B䉻%b���F�s=~)����.��B��*{Nd��jI?a�>���`� #>�B��L�r�c"�,lf�{�i#r�B�)� ��1�ɴu;�%��<O�����"O��Cb-Ŕ[�di�+ӤRy�$"O4�DkȆU�e������;�!&D��wċ��� ��!�"Q����v9D�dCg%:"N҈{���@�~���6D��h��V���f(F7�f�Ceo4D��S����@d���Ƈd��*d7D���Q
�5�Xy�\	�e��)�>�yĩ�8!��/��q�4)c���yb�_Ì,���7<�x���W�y�gɞf���臂X�4D�[#�K��y��A�Qy�-h�02���#�	���yr@I*aߢ�0�U�r��� �J@�yC�ad�qg#��k��%�w�Y�?����}�L8�:p�\��QFv�&Y�ȓe&���si�)���zw���46�ч�e2��e���Ce�N40�00[v"O�I���
&.���Ig!� I��|�e"OV����Q=B4HP���@5"O���C� �����ƗXe|�q"OZ=���H�M)\XI�@+\�E�D"O6����ugh�Ȇ%C�d\�"OR���?a��=�Ec�/l0�d�"O��5�^6~H�b�"TFJ�1�"OV�	"��%+�A �� b3�X�"O��7fS8Gh6�QdW�#
�h "OH��Ү��h�~Db$P�Ƅ
�"O�"䤐�G�*]8�#όJg
�!"O%�C��f�`�H�"�lI�U�"O����͏eB8 �ŀ
7B��"O�y;�KC�2}��+�/�2 �4"Obej�	`�)��;�؝[
�'��%`�nA��pA���P\��' �A�(7�NA[�"�	M�x�'��0�m:c�l@�aE	6�Eb�'�jh�̂;a�nL�֩ ��<`�'G$#���[����Oۜ�3�'������b���a���@�'�����	'g@�3�`Q2�z�2�'qrXh!m�:QBa��(Q8/�1�'� �b� M�p�+UO�����'��ls��;J�A&�S�!:�'�p��m�{hD�@�����9��'��ɠQ���(����`�#f���'������/6Ժp
�"oت���'�8y� a��#^8p�sD��x���'�r�٣�=
�&$�'�E�_[��r�'�\a!��ЂU�e��P��I��'K�I3¯�5���s���Me&0��'I�����ȤO%c�̚�s�d��'�(0i��pd���͖xL��Q	�'�Ё��fՆ&���2�]n���(
�'F��FJϯ,����i�:ha���	�'��Y��hϚ����3t�Xe��'�TIC��ŭ�qJ��=zBe��'1Č���;l��ĩ�lH�:�$h�'�� IKE�D����UN����)R�':�@&�X�aʰ< n�b���'�6i���*@C��U�ܹ7�tC
�'}j �עT�K!*�I��N<(?P� �'w�c���3̤Thu�IM1��
�'Kl����:��$ĆN'X̲q3�'�T�	��^6W��q,2�����'�љ�AN5.
��a�/m~x��� 2|ra������35l�S�v� "O� cv��+JX�M�W� �C�"O��!F�ߛN���4��&R���"O(K�l�)/̃���+3\yir"O�������,x�J�%h�(�"O��&�*���c�[7<�F�:&"O>�s�i�!~x����M(J��)�"O^���A/,����R�F����"O�a�#&ی��9�Q�N�Az��W"O�e�-]�c�`�5�'8��\ �"O<1p���4��7�ġ�<ى@"O� [BO܎;\�<!�]xw@���"O��"��	s�����1T��k�"O$��'ۧe'�@r扝�ND"E�"O���ЬD�t�=��cQ/{�d	ò"O��1��%}x�@Cҟ&�.cQ"O�I ��9�����է;��,��"OXa�P��_J(Ɂ�F*o��iz$"O*��O�r�)�:`���K,:!�$ۊ���"��]46�h�U!B'�!�D_
(�����u���#�f�1!�$C�H���'j���#$�a��B�I8,~��ie��fF6uh�c��j��B�	=C>$!�c�I%D�М��B�K��B�I�=<����U�*7�4���3tU&C�ɨXP�1X�!eav09����J��B䉙?�\�
�"�+�L��5��<lY�B�	���ը��-��p��KkB�I��f-9���"��uaЮ5E��C�	�1~ޝ@�L�Egx"�G���xC�	�.UTP��_ tt�B�SPC䉙U� -�b��-|�$�:W�	�.C�ɋ1�,x+$�Q.�
T��a��B�
Bcj�����Q��I �E�G��B�	�\��E��#b��}��JĤ<�B䉼/}hIx'�O�p�w�±wlB��{4h��\�<LK7m51�*$"O~�/\q��8{�lW�)ԲUp�"O�@a��JL�pW�R�)T"O6�+c�V�\�c���	셣�"O	�!	�<�Wć
�P��"O�h�ӁT�:-�l�b�!� �3"O�x��E].C��V�-Kz�T"O@1����2oh�Qd�OFbQj�"O��_�"�����LG�pM� ��"O8�q�G 
-�������/Dxe#"O��QF�S.5���Dj�+4��P"O���
��#�Р�Ș�'���"O:|�4�#�d!��眔	gr�j"O.T����'-���TG_�U�,��0"Odq� �@��!��

qI"Ob���+�7Xcv@��% �d�n��"OPb *HT<r�ß�WQ�"O�ݸ�I�V�Q�(J*��"$"Op���-�߼�eM��	BT��"O��z�>�Ԭ2�!6G�`�Q"O^DY�D��=eH��ǜ�i���a"O��SJ.FF0��揜Y����"O��e��:"� LH$��)N��%��"O|esbj_�M�`$ƪ�V=2�"O��*g�Sd�p	�wR!1����"O|t����7��1��aӂG��A��"O��9��Xh�`�;�M�{�ṟ�"OJ0� �xذd�֯Ҝ��9
"O� �J�g�I~�m��5y��
"OZY��d� 2�Rx�K�]pj�$"O�X���Q$_��ز`S)XU(9[�"O�y
௉�+���ЅXUx���"OHu��9xppHӲ��-:*{p"O�����?.u�����k>U�@"O�0�D�:A�X�1O��Y:��@"OF�W��i�8��m<l��1'"ON��u�� 8f���0#�@��0"O�TA��h��$
#�9�*��"O��UA�}�ʌ+�@�^��9j�"OҭÀD�o�QG�T�7�2��r"O�y�ń��`���	V����W"Ox���hK�qn+hb���&"O$�Se��(.������/X�^(��"O&�8�� RabL[���-Q����"O���!R�y�D������2"O  8!�T'Vy��kFU�:0�r"O޸*q�=D�����A,�<��"O�`
���4D�
6�̈3���G"O��c�לX��A���C)�x��"O�d�fCz"r�	T	�D!�D"OZ��'b���Xs��%
�"}�#"O=z�*8.ڸ����4�X4"Ojp���E<S��LyE�N�C �9�"O�	���/a�����ڤ(造[7"O���#P	
��D���G"OM��,B%$. �84 ĂK�4jf"O�xLM�ʉ���ف�HY:g"O$嘔��u�nAXԎD�-����"O�Q��5d`N� �N��]�\�"O�*=��:�MQ6�v�ӳ"O&���d�'�bl�w�@�9uMcG"O���)�!�S��q>��1$"O\!��^P:(E��R7M�t�"Ov���C�5U�����W� ��=��"Ov���ժ)�����Ҍ��5��"O�uQf�P�A�&CB��,_
d� "O��r�S5C����a��s�Hs�*O:���	i}�,�b�ّi���	�'��U����[��K�Ֆ-怔J�'V�%u%]�0�MH ���0��'�\�`�̺�`���	Y�F0)z�'Ĩɤ�	��R��(4GPa��'i��%J
�4�������p��'ߒ�1�d=�M�W�:i��P�'��͂�F6n5 �dMc����'�����\D��p�hԶ$($��'�`���	Ί{Ȉ���_.4��@
�'t�%j��Ak~3�,�c+D��' D=�A'�&� ��
�e��DB�'Qnl�t�<mja0��[ZP�	�'�<}��b�kH�l"QcY��i��'btp5��%Z�"�)���>�����'��,X�T�L�jD�g�F���(	�'�U�CF
ul�;pa��J�Ҵ1�''� BK@*7� c�m�2P��!��'��xHP��.m~ƨ��۷W�5��'�"��EW"V�;ƧѸV�t��'4
�h�6/�<R��ɯM��8��'�P8���Vm�����F���2�'v4�#vD���D��A��9��A�'W�q0�*��,'�����'$�tЦ���\�T���m��.�T�B��� t\AGZy���Q B]\��25"Op9H6
՗���v��I����"O0Ph"�
G��3��G�2���3�"O�\�u�H"u<��YO�7 �r�K'"O:�X�e�0G9p!����x�2"O��"�LZ!6�`�w�ЖI�x��"O���c H�y�kD�t܆��"OJy(3n֦	�c5)H5x�<pYQ"OhM�U'��#�VD��mR��r�°"O��cé̳;�"P��(.�Vȡ�"O
%��	

��sc�_/P,jb"O�1qR
��q (�7y���e"OZ�sEdO ��A���Ϻ`T����"Oh���ů2��������*��"O��9�NQ��6��F�
#����
O�6�S2��
�]�Bt�
��?O!���ޢ��X�uRqc��D�O>a��O��y`l̫{6T�Te�w�,���"O�My�����d��F3g&���'��,���W�^;!N:/�����f��C�	._Z�g�	!	1�PCG�T_�f�<9��T>U8e䕬*.���
� 1�G�?�O4�G�Z�Jdf\��8��&@�QnNAp�>y�H��DD��'���*u��C�4��0�T�)Ū03���O�&PG��KN"Wf����
���s3.�	�����D,����'�ȅ!7��L�*Г��ɪQ�� jx�J��?%>1+N>�w	Ӏl�xhŦڤ	���X�C@T���=	4Ą�4�pti��H�H��z3�EO?	�4���`����O��X��I	>c1���������	�'w��횾^O�����@*�U����'&�>��5|��x�GL�m�f�N�s��B�I�y%��7K6���rӾ	D���K�Bܻw"�O&�����6`{��,]P� pO@�=��p!�"�� ��-�ȓU���a�L�(�HE��ӡih�8�ȓ3}���m���0�[2��}�ȓN�:<X��YFT����/��'-a~"��;v\���m[��r\yvm�
�y�Φ6����� ���ɲ�W��yҪ��#�@�d�o�|5#���y2�LY��"6l��a�*{�&���yB�	5p�q J^8��zC�O��ybd�B�@���\T.��f?�y��@40��3�_,Z�Z��An[��yrb+[�\����߀Xh|T����y⭀)�@�8�AS��H�sꂚ�y�F�9�#�s�:q�s��ybϘ;߲8xtCJ�V�й�!���yr�$ �DTPn
�!��v�1�yB��:w=�|!w�ߨi�z���]/�yBD��^D̹[G��U&X#�����y2�]q�����/T�����G���y2�݅0ʨ�y���"��|	d�K�0<��D<Wz�<K�/�(@&��	�O!�đ��<�{AjR�,$�2���j������j����Jn<�� �B%"2*S"O���*�1bT�)rUNġ:"�|˕�x��'�ܩ�J��z�(!�Nӥ����'Q��� %�E�1��=���'2�p��$�	?��\"�b\�9X��'R���g��Ft���jەu��[���d> |܋g
U�[�,ѳe-� ft��r����)q���vdx@�"5e�yӧ��x�O�I3f$�`��9%�Ԋ`�L���� v��e��p�� (�CX�~���v�xB�)�s��9*�Ѿ3%� �%ɤ�����>yy׭'A�v�"�V�N������"��[��V /$H1�d/D�t�����h``-#h|�sO*}�f?���'q ����9n�ޡ�@oN�7ƽ�	�'�p݈#��~�xS��+x�lA�'��|�e��a�hp �0Vb�'�铎hO��5	kn��f��u@� �B�z����5}��6,�ӱ�$J��11	�(0=�I�<)览��
R�ʕ��A#O~��q�ͧf^ay���O�U�c�=F�Ь�7&&$2�\���Or��M3˓f�<�8c擿f *	�u�ў6����Iæ��'��~��	!��o	��o�(@<� �$�2D���"���V,`�f��,ڄ
FD0��8�	C�O�|�X��tq����P�X�����'�(�X���o㈰@�hQE��M�艈���ʴ~�6P�� ګktj$X�	8��{ң�P�IQ�^���	}�ƐX��@$i�Tc�l��I|k�1pAf�
R׬�3��}Rb�L��~�;O�'�y���KUR�3𤎘&�0��f��y�o�+��� �˴��44������Ly��|Zwn1O��)�>���K'C�lH́�"O�|��K�;�}�t�M�tjt���'��O����ԟ�(J�Nѐc��A��&n\֜ �"O�b҂5�@e¦��7j���'UDy��)�`	��΄�&i�p�'��D�2B�� 2��@HrA]W�\S0N��ʓ{Ij��D.1b����C	a=��QnD*M�1O�=9�'��IV�>|��hK�t��Uꛏ.�B�ryni-�,l�Aiؘhn����-�'��"=��I;���jV]��Y��ܥxݤɇ�ɛ�� eH�RSf]!'�][�bR�^(��d֫��'��#}�'[F�J׭)��)���>�Z$h�'�����M#t��@0�%�#��Dp޴��d+�O��˂��7
�I�(Bo*n�s��IM��Ҧ�()��j��JtMC��l��Y�P"O���)O�i� %C�G�l�p����V��?uP��[�X��W��5W_M��C3D����Jp� �G�B�`�@�;D��eE6]֌��7�2+�����=D�$�4�+_Y��J ��7 �� W�6D�`
�J��_�<)�Q��`���K�0D�HPc��:q*���"� 8�DБ�J0D��q!�6�婓�حZ�"l��;D�L�%N��C9h�+"j��ռ�h�$;�O�ʓ59��r��^�>i��_+[�~)��6A��* B���9[�<�NĆȓZ���O��
��j�$h���`jb5Q`n؇YLrt`�&��G����O�=��&h��dłdc�G��|���w�<�G��j� 4�c��=��}��ƁK�<�mK�n�V$B���(<��,��RG��|�?1uE�����$#�!���x��A}��'�� ��W	
�xk�*V>
3*�B��~��'�����E&e�\!+%!¶O���'�|�J��Iz0i���G�@�r(+�"�)�4lb{h	��(�%k�&5�S��yBjX�Qz|	R�ΉhY�쳷�A�yB��B�֭
�a�S�N�j��Y��0>!N��+��88=�Sd�9Kg��C�K���+�O^<���sc�c�m֝Z�h�s2�'�qO~�D�\������9�@	�NO6!��¿aOЀ��މD��e�,=$�ax��)� 
q�@��@�"A��U��0)�"O )rS�>� �h��"���"O��@QDD�x����H��x�"Oڹ���N4�nQ'��:P��4"Ot8T��7vf|��!�Sp�	b�O���� Eވ�F-cb΄r���	�'jx���cM�~1�l��DG![����N�(�O�=�'4��Ma���$���Q�U��fD����{�	9W":�D�̬Ws�Ts��R0r|�b����	<"�)�ܢo�.8����b������\�B�t�t��� $:U��$,?1�(���j`��b��X����N#z��ȓOpDh�+�B:�qx��K
0ZN��:�Hz�̧f�x�`�˞ �e��t���⚔�D��#�3���ȓ7�d���5/�xuÚ1�ڝ����u0q��1��IBp�D,{�LP�ȓ6;�H��n���J$���J*
O���ȓGE�AC�J(S�z�y��P%R@8���D)�ݡ��1���2CX:R�ԇȓJ��|����D٤=��O�#�
<�ȓ%���)�NHH��-�QM��]��)�ʓO��
��ş\�^$+���)`^�C�ɍ!�T	WC��;�@��u�_K�C��)7<�t�O�7�lq ��"o�C�ɔX���Zqg&>
�8����y.�C�I}��I`t��^ �Ӫ5}?0B�	6�����6P�*\�B�w�C�,��d�� O7g
�`Bc�oj�C䉻 7�2w�b�c ��C�I�_�R���b�7F���N]�-��C�<| Ea5Fَꆵ�æ\��C�Ɉ2��E�ԋ��"�()�R��.X��B䉫O�H� WAB;z�\T�K�qA�B䉨wY`2$���6�d�0��
�KI�B�ɕhM(I�vd �N�`` �I?,�B�	��0j�D�6[�BH ��::C�Ixe�1*���h�� ��`�`D�B�	�-����J��M�@b煓��B�)Tmp%�P��8B��|�S��>H�C�	�K&,�Q�Ԗ��t�r�ۚ|C�IH� ��0"�;!،��Z�"/�C�I�%\����w�n������8�C䉦244�a�eY;9y�$+A*��l�nC��2N�Fs���6��P&$p�B�56.�Ms4��E�AI�TB�ɕB�1���.uv���Nҧ�B�ɀK�-���qGx(���K2E��b��# ��B��0�TA�fR�c�d&�ɦ
�@8#��՗e�A�g����B��c�B�{��
>VV�0��dvB�I�{!�I6��8�"��@/��B䉗k�>����
`� ��L�nB䉆>�&��1�I�Wؕ��eN�!3vB� OR��N�H@��a��mC䉥�j�0%�S ¸��<�LC�	l{1s��ձB�*��\.J�
C�	�$׎�x��˂b,pEq���6��B�	�iv�5P���a�\�� K�B�ɳ*�!�u	;nQ��AdS�)m�B�,3	:�[� S���e�u�LB�	�x&8"�I��T�p�H�fN�t�B�	g؀iQe�F]k|Hȓ��N,C�	�ܒ ��2b�^4a��9V�~C�4��䲖!�/�f��'E5s�rC�)� ూ����Hmr3늁U޸!w"O�K�D ����d�0��@�"O�ժ0a�OM&�ƁO�>|LU"O�h���u춉)�.�U�4a:d"O|ĻA�Ј�u��n�w�ry��"OD�B�/U��iS�CX)�>xg"O��MĞYev��!�߾6��DQ�"OB`c�N�/}H�h�E�څ/��=ҥ"O�ͫ��G�	��-�x>� "O��؄�Q25�w�ֈ]{�8�"O3sFĹsdN	q�J��f	<���"O$��f�Կh ��z��Ϩ?�dY��"O���dŝM��@WF�-�0d�a"O��@����_qrȪ&/ے|l�j'"OB� �oU�&�
IHDϐ�kz����"O�l�¡ڋⲁ����ҕ)5"OD�$��n}���	b�BPs�"O�����6A����*#�L�h4"O`�IP⎋mÊRnA�t�)�0"O ��b��h� iۥn%�h3�"OF%�7hТ-Q�d��@���J���"O�����I]�}yvl�E�B
e�i<hZ�'4vE��l�5d��y�'L�O}�0B�w[b�1�3?9�e�;�TSR�Z�N���Y�#No�<��Ի^�r�딓Of�JC��Nܓ2a�q2''�����9�Ɯb��W�&�nd�B"O��a�-	�x��U�Z�s��ΣrqOƥ��Y�|9��F!_��+�l�-<�ܨ2D�����L+�� (�|�X���M\ʘ����9�O��L�9%�pT�B�W ^r}���'��e WC~R�ɂ"�x�#î
?�μ����y����~H��AD��-HRƌ���'	��)C���ԍFwh������,;��@o���y���%kA�0��9*���y��S�\4�t�͔{�"��$���y��!E<����(&��iy����y�`_�s�-�� Be�Y�c8�y2�3xUd32��T��ݹ�ybHʶ[~�!*���4(��k�"�y�I��Yci*�O�/bz�Zb���yB�0o����!��q�f�ڦk��y�
�u6xup�J�t�`9S!���y"(٣h��`Ѫ��bKj���(���yr�Vnbl���
[2�q��K�*�yr	�dt��DQ�On�4�c���y�ǎ-jXD�Ə?@���B�L0�y�N!l1d���!lp��� �y���^��S��}��1��B�y���3�lHc/߹r���s�A���y�LN9<��I��!��`��I3�$E��yb�^�*8�z풛������!�y��d�f�0ch�JP�DN�,�y��L+-�(]R��4<�$�D@L��y"'���{��+ \��d& �yr�0L%<T��2W֮�����y��^�A1tP*;�`4���y�*�-P�M��5�����-��~2(�Q����O ������=���B�,,�Wt��wj߆F(V����Q�< b���OZ��c�����%Oۂ���:O�[0�� }�O?��%!��hK;b>���eJ/�	�=�@�iU�!95,�!��])2��ҥ^lR�I匝Bn�	�ct�qq��2wsay�CB"\!��r&��F�� ��텸+:(���
=(c؝@D�J�<����[
u_h`䫈�:� |K�KM�|h��)�
����ē��8#�&:Q��m)���\�Jm�	�`j��sŉ�A�P����&	�� kf&˸U����� >a�-�f��	R�'��dG�q���'| �D$y.ICGm��y��Tp���3`|e�`��5tO�A��)�B�r�hsf�f��3ڧNʖI��䇓x��D"�k�/Lv	����/d?����!�t��d��$��ĉ竇�=�!���#J�	/��kDl��z�ay��[
(������j��,��J��В]�_����v��?I��D'(#�Ua���+F�@j&��L�Zȱp 
9�q��I�y��Q�Q�,d�Q VI�� הt1���tq�fڄa��[��HfXb4PG`�6.f�Y6�>a�O� �Y�n�;9���f䔞%�T�����N�vV��y� ״#��8�����k��H��ϫ3��ih�e�hW�E��K]�1��2cm�dZ��6�ڄ��y	�S�$K:��&֠q�C �K���q�Z,��˟ �pD�Eg�{�xh�Ќ��iֶ��L���I�dq�Lc�΀v޸|�hE�-�F :q
ɉt-�@��'�R���*D`��|
�EY��>]S4�>z���Z���>A�iZ#1���c��V3������0A�ҽ~��i��	�g�/a���,C�Ne�&,��}G�~��=��<�s�[�IiJ�����H���Î<0��oZ4��-�� R�6��S�b`�1��%�Z({稖�-�f���j[>�*�D}�	E�r�t��b��[�'W�� ��:f:�P �	�\�FeHŘ�x� �i����H|�>!�a��J�:X�t�Jp�X�I5
m?��!�UYZ�Ô�/}��$%�����qa�(.`��A��hU���@Ω�Y�
��G�����	'E��Z��l���Obj5�Ի8$�d���"�>-��� T��'G@u�Q�DFa@�����::l�˦�'ƶ=3�m��G$��T͒$]! l�S���=��5K"��<�%� �<q���<E�t#)z��ȃ���w�*͈7Ğ���OJ�c��^l4��>5X���([�:�iS��<N��A�G�?D�H�#(Y��z�jU�n*����`�<���T���OH��՘O���v��5�r|2�i_�Jڨ��'��8�D� �1at�ж:B*)z�OC�H��ow��O>�˒钼.Z�q��L0"�� 
tA;D�����{$蜋�L�&�t|cҋ����,WH����dWl�3�ɭm�RM�bnÌxx�8�'hC�(�N���Ԭn�F	r��Ƥi���h����O��铩"%b\���>a����]A�
A���� ��ER$�sy�ztES��3p6���jp��)\�0�R�A��6�3�N�un����'bH���LY,}K\:!Ԝ`�HYy(O�9I�hՇVy�q3%E����4��V�DU ugv�T
��Ɛb1l�2T�����ܷ�y¹��΅�)����A`ת1�)��eJ�{�P<�"l�?n�B��"OZ�>�:��ݶ�yWG�/-������1pV�Q	Ǌ����?���*Wpe���*~ �Ѹ��CX�lp��'F�S��G�r���.�"�*���4�D"�̑�ݤ�cuʘ�$5:�?u(̳Di@l�&oU+eB���dM�4P&|���Ť#�쥙vC�7d��b��B^VFd"�>�O����p7<]�F2��T�W��|���f-h�&/�2$[��:��&Ht��(&����	H�����чW�LG��P�Jӣ�!�J&ATN(�!D�J��B�)�xкDB�eš'N �da�, ������?-�BĠK��RҩK�{��|nF(���=K�x̺�BUv�a|�#�4�0�+F��>5t^Ȱ �#�r�C'M�G�V��gԃҨh2l9w�,i���[qR� `-�;?*=�#�M"~�:WҲT����?Q�jQ28qpLR �F�8���&`��G��� ��8�\�q��R��B��y?�Ȩ��5OLUH$k�kuB�;��\���"~�<�@��U/����̔a*65����(�=;�B�/9��X�4G��qR_w��.�@���Ů���$'��^5�������C�>�r(�/B�u�mZ� ӊ-cㅒ�@�~��ҤZ�A۰zr-X25Y"AK�mV.@�iH4�[�%Ԁ!C�e��E�󤇱?WH�@�=d��L���N�����F��=���,D2���-���i�-��H��$��8��<�'iU�`�V��Ä+\FVE�C�J x�B�06�Ŭ��<I".^�`�0k�(	(P)P�a}���B�H�x����#*q���S���@	����Y�⑓s�Tl�$��HP��qD��K���3�F8�;ׯ��?��W��xJ1����<�yMa�Z�	){K,��PΞ�[���` ݚ��GD�
�u�!�8�x 6＝���W��АG/{��1`�	�!�@I�����6P_���?G���BJ�Vd(��K�b����(/�� �� �1�.��NW�E���2����n,H����L�z��fNZ�>��	�N�ȌFx�	[�V��y���$mr���)_Q���ͺ�D�S�A�D��\�@��)h�̄��O?v�(X�<�=Z���)������ �]o.��'���r�g�|���B�6F���AJ�)qwnx� VH+�lo�"|iT��E�4�}��'J4$B�ɌV�< ؑf�|u�(2a�4}�*�x�O�QDb�n�
a�a��8��G ���O�ļ���JM� %/D�a��M���|��̳�%�J�.	S3∇xb�8�卓A�����R�1(�t�戓Z�0e� d
�I�"C#R?c���/�8
;Є�׉�.	���Zte'O�Y�ц��L�t����	� ��yU%�����s�釐p8�а�aKTR�	a0��E�|��	�<R�됃����gJ�& ~$�'�B��vy�$�f�����R�<�39�j�	�ˆ�dn.��F"5PR�	�"O�E��vB�@���	Ul���&�'���yGdM&l"��(u掏o��A� l$]K��d�@^����bƜ�V��� ���=y�AJ >���OLp� 
H�>و&ϕ8YҠ"�w�$ğ.$d�$���С��]hԍ�2�eqv��qO�0��ʃ� �d�"�@�pD�ɋ�v��I)��9i~�"�� �s���@��'���C���&x�B�n��D��5�T�=Q�-Q�<��ds>�v䉞F�ֹ'�L����?A$2� �C�(
���3D���M�/lp�� Z�:x�3P��j���a�q&��$�b�1� 4>s	s��@@�N���I�@�ȀKP�Q�/�xnz���N�/Q�8��#j?g#���ȓo�h��V�yQfD�D)π����=�ć�
x@ZL����H��ݻ�R3�z���	K"y�}Zg"O��H7�Ͻ_� #����N�qi����m@Ay"��y���6*
|s	�58�퉱��!��@�:�a�eL�� ���[4Y� [�@�u_�8;a�Ap؞�T��-�}��,
7��a��&lO�Ma�F� ):����f(
q�j�lb��5b��@HT���m
�{��UX��Ibd�-*�&T�?�e%T������G�_�x�NޫAn`!���n!�D�=0hd���)X�c��ƶ,�!�$P�t@�q�o�'2�ݹwg�4�!��6=�4 �r��	~]`
�,\�!�D�0^�>��&I=S8�E`�o��W%!�G�i*��2�ߎ/�P��Ł( !�d���D9Q��t�B��p!�A�B	�%�6�̔`R�9�×	g!�D�	!G�9��U�XP�����M�A�!��]�$H(�l�)V|���ѣ�!�$B�r�!JPo/Ӝ	����>�!�d��1��:c�}����`��6,�!�D� ���C�N�s���`����!�d����:����o�u:Ao�>e�!��ķw"�P��� !�4A�N
�y�!�dK�F�>$�g�]=�T͟�Ob!��U_88`C�� 'R>hPN!xS!�$�o�2`G �
'�����S!�d$0fe��a�} �P��oM!��J.{O2@P�Ԧ�9���D�	[h<I"e�oJ��ӥ�8yR�F��I�<��I��b�@���ۇ%$�!��|�<)��Y� x`��2�	=�$aR'�}�<�A儦Ǯ�$n�?s���h�KH{�<��,�*{�TM�&U,�L{C��H�<9��%j��`I�!�<C�m�\�<q��E�?Xr���IL�.�8��4BOB�<���@z� ����B�@A[�<�P��5>�Kp��{��r�GSU�<��bN*e����7Ď�{�^�q��d�<�7F�"�*����dbbA!�d�<	��f�������x�<q��Y��
	9D(߅�V�s�]R�<1'μc�ֱ#R�"����*J�<�CFƨ���,��<H�A{�@�}�<�L�0*��1�#Hr$+5i�x�<�e�S�fx��q���(fPmf <D��kŏɬr�u+dK�,x$���N1D�����%[KnQ �u>0�Z�$(D�<� �ѕh�^m�n2G����;D�ԪE�T	b��$�'��2?f�aj6D�iw���%$� �)��D9�}
	+D�4�j�Nք�B7(��L��X`�?D�� h�!C��5���XvMA�wo mc�"O2�2�ȅ�-�!�gBE���}�v"Oda�H�8)m�y�dA	�g���"O6dB���>'tf��Vծ$���"O E����~y|5�Ǝ��c�P� �"OJ�
��,+4����E����r�"O$��"�ة�Mb$q�����"OjŰ��^�6�b]��d9�JT��"O\Y""k(��ᢱ�SBu��� "O�`Hb�Ĺm�=Y��P�hl���"Opl+Qd�~ͨ��'	>C�ִ	�"O�����e`�f�:Q`$�"OL�Q�Z�\&u+�(��2Y.e�4"OH�y	E<�!1%�:qGFp�"O�aiQ%_�Qƨ�P�В:",��"O�t*gŔ�m��i��!,z�!@"O,T��(+N���5g�4,\MA"O����0.��Lң'�� Np#"O< 4n�Uۂ�s�]Q&����"O�<���2,�8I�E�4�x��v"OzѸ2NQ�)���0�߯f��Z!"Oƹ:�NGe��(�%�TL�u"O��p��CN-�c���tw��P�"Ob$!A��1�0@������W"O��H�K%�D��84�L��"O��0��\<z���FSC��h��"O@I#pn��||���M=Rxp`"O��҅|r��6�˦Z^���3"O
9Z��$M�4�)2$yS2lrS"O�-���Z�@��˛h��ps"ǪR�|uLM!�ꖪN2� �"OB`�"
>^/HTp��uC���0D����G��us�S7-$V�[��5D�1�'�$5�����4^$ �-0D�d�V�V�޸��_���	b�/D����BOw�ĠCA� V��I"�,*D� h��ķZÄc���Z��i�r�6D�d���C��hxek��*�)YL D�t�� �"Yl��"Q,J8���bI-D��QpMG<��@���+w,x	3W�-D�̘�g� &�Ys �\D3V	(D��Ô�O�.���˜�~�E�A�)D�\y� 'fE�3E�B�Yh�n%D��!#� <����S��BC���.D��÷�"`N��sϘ�E�`��.D�8��d���a*А�|At�!D���uO�tG�� qK�l;,��V*D��1����}�P���t����<D�)p!�30դ8���H"x�2�3@�(D��	��Сgƪ��4䍏x��A�F'D�!��:u)8�Ƌ2^-��"�G$D���ph�b�@�V�.���� �#D�da�Ǚ�N�y�Wc=|N�$[�o D���p����8C4�I�Y�^�+E�*D��[ueĩD�
1�YHW�y� �7D��	U�8H4K([��
���1D�hB�m^={$�i�"\+��l#S�0D���D��:�qT�\�V��4�p�+D�X2�n�;Y� ,�)t�x��`=D�H���T;n����CG�TL�0�>D�����/�u�f$�x`6X9gn��x�V�5"��*�މ��0��R�P�l�<} �tSt��p�P�'����&��k���f�(��A֛=DT��Um��y�Ȓ�n��S�|��)L.#�qYŢM�VTɛc��m��O.8����_L������π ��ۓ
R�f?��eͱE��t��\��P$�6����'����]�vؒ�k�8��F�I-**Q���Ǭk?dT̓��O�"i �M�ZX(a�u�%����L��K��с�FH<1%�ʕQlh�sp큺(ޖp���K�T1��G<�
�����&���U�KUgh�;��>a�OߚQz���N�f�Xa"��vE���ߓ#|��D�_׎y*#n[$
d���&J�9�d�v)�9� a�%�U��4:�`�'�>Y�w'ƾ3dd��Eg �ڠRW�Vs�U�D�
�o�~m���Uk���O7�=�բL���p�._ Cj��-Onr�CԸz�z�	˓*ݨ<�&E�@K�UZ�b���䊲�KhX@hYtdZ�/,���n�';�Q�����rݢ⛌0�P�Z�ڹ�d���l7�O�5/L����E�:��d�'M�A����B�x�M��MP�hD��)y��9���D�>��L���'yp$|�-'*��)2�A:f���F~2���,�b)A�l�p�%+��>=��ۀN���a�L��O�ոrN���<�1aX7_Ĵ`ل�*�"���|�|bK�0;zt �����+\ 0�q��~�C��wZB@�R�I�#����&�>=�`y���U�dMM�2ě�� ;^X��x��¯6�h��̜�<Y �˥�'(�z��F��\�Ӂ�p�����Io�|0�>ƍO�fO�XS���b���aH�u˲��0��k�i�z���.~���%��m@�����)�O�aK�hD�E?h�P����Q��Y�$f�3��$(QcF�M�B�����H��f�]~�O��d�R��\}��ťd�r<
�JT9O=�|IC��٨O^Hrv��F�J���d��&v���:C6�SBᚶQ�(�t�x���h����'�D��2�J�C�0!ғ���i\Ԡc�'T� 
F���	�E�Oq�ԥ��JM�
 xu ��V	�|�6ɀw��������R�a��:7�ji��7�|�1,԰��$h  ��c٩c�ƙ�n'$x�F"�č�H��]*g�3j������;}�2��d�0�,�feU�b��!��Ѽu��3��IP\ �'<�Ca�9��,��[8E`�T��DQ�fʽ����(,��=*c�d�'S#��//�䂗
�61���#�I-D�,P�O�6��9�n"��˒��<ѣ�����O�����Obj��T"�b!���'���~
�'�*�
�C�1��e�ea]*�����O*��@k��VF�O>�t�S�6|�-�����^etA�V#D��!��%Ű٫'&�2��x�#���		`���p�C�3�	�&rt�a�K�Tɨ4�Y*����%z���oR��^Հ��N$��8�8Y�*�X	�{[ʽ�g=U�8��%d&؄D�n��Ly;����N��p2����ՅQ�8�� �*R����x���\_���'��A
 �L�[�,��e�0't��-Oji���W�HrΈ��W%`����7J4j���G�I�4�O*�Z)�DƖ"�f��"���yҩ���l9�5�H?n�f�ejR�s����`)�_ъ��v-�;U�0�)��+���t�T}�>�Q����I¼�ʡ��Ɖ�T�'ǾI�a�+���y$�-��=K�D��V����!%�L���Y*$���"tK��VA�"=��dN�u��P�� �7o�ANi�'�1C3��{ڶ%@�d=��4�� ��3��YpkP�N�.ݹw�2���k�b�m��	7^�1q3����f�@@(5�"�9���a �Rm�uz#�
�$lf�����/�*�V?FF�:+v-��H�%�y*U�>D���R�NV ���J�5ԚuB"F�;-��t�Ńڮ�k�m�$#j�����NR(���J:5֞}Rhޅ��$ޠ)�d�I�_iF%��)�OH�jc��'BN��O�n^��å:e ��� [�̩�吋?V��fBA��)I�O\�Dz�m��,B(��aN�~��W`[s�'�x[�e7r\��~��+'�۲,޴��2*#�u; �M�p��1J��;$�X"��6`������`Z�)͌b�d�d��N`�A��a����'��d
�y��&F�t7�"C���������1Rp�H�DV�R!�C�Il|��1��
D6��2iY	h�P����ߦAIhǾY(93!�KU���?R���''��O>|.ufՔK�j�����u�h؆�ɏ2��HR�={N\�[�#���M���ѐU��dR� ���o�o�<����85� ��S��ۣ��Gy !`Bm��O0�;G�MC�O3�ei�[�%�T]X��G����'Z��b�h*?�x����7��[�E,�r�� �*��P���gܓ naQw�]��, ���,���	?"iQ��Ãt����=]��u�ʉ�n4(ig���b^���E�'}��AS���5���W텟i�*��D�X�.� Z�@k�Go�����/X��"g�L*��b��y� C�I@�@!��u�8l[�
�LF�Iq؉�p휡+�6)�F�:���n1 ���+H��@�N�bX� �'"O� 9��Q{&�1���[괜y�s�$Z>n��Ais�1���6w	�d�ĊX�z�l�.�3&[���G7tl�����L�4;V���X�(�s)m����?i���H�c]1+��{$(�����D�*xQ�=����!Z�Tl��W�!�!��_*e��/��sk��j4k �6��=�����H6�)�S�o�b�*Y���+�B^_��C�I"f�P!	3�]%0˪��2��8OC��$��1��]��:�O���%�-X�&��W��u�H��R�����BkՖ�d��<
�bt����8�⤇s�!�č,<�6족Y�g�R�a��#�qO�!o^ij��A/�'H����3$�)�e�Y��[T�R�<I��Y$���0�b�?��3����@P�]k�A+�I:8�Q>�v�<��)��2�r!�6�	3R9��yU>q�H�0h6b `�
	+��%�wE�K��9�cǃ�a{���8H(j<�/�)�r�aD�P)�p=Y�
�Z~ mJ�*]��M$*]���q�uc$nMN�i�aZo�<�4�U�p�~AӡHK +�a���mܓx߾�h�D��D�#��iP��T��I�!uf��0�Ӵ�!򄌽+X����^g)B�(
���"���Y9�i�'r�0D�,O܄0�ԻVz`��2(�p"ODt���d_��.K64�K'p�`0x��Q<��%�퉔	Q��� F�^���p��9��$3(����ǃ�?A�H�#'PP�/�"7�.H���v�<	�dE�L1ŋ+�Lyґ�O��O8v��1�I
������hWD5��c�N�1jb�*t"O.��6$ZrƲ�Y�l�=���3�"OX��vi�(L8@:PJEhO0�c"O��eg7/�v}rVh��,: ��"O�U��(�+�I��Z2.�}��"Op�8�!�,1��Df��-\	zG"O��Y�bCO~�s	Q�RDK�"O���!+Nn
�c���.!�݊�"O�Ƞ0����`�/�*T����"O&�:� �/W&8��/�m�:��"OH9�"�FQ��Q�Q�Ȕɠ���"O���E˺g�X A`�R�G���"OnTXV���'y.������q;�=Q�"Ob��gMۘmf"���
(U��qq"O��-7��<2 a4(z��"O���'枋U;B�i��� N2t�q*Ox{r�W�#`��:�&�{x.��
�'���"!�	���D���r��Y�'�>Q@��8+����ɜ���'2 ����ˆT1 �8�&ˮF()��'�@̋1fF�nk��"P��j����'����"a��V}�H�p�m���K�'�-�ɕ�4���KS�-S�(�;�'\^�9r���J֙��#]�|@ 8�'TZ��V����U�ѩ�w+4�z�')&�P24�MhP���dt�9�'4��s@ݥ7�\�'�U�SnP�'�lL"qa�bV��gքqd�p��'�ԚpE
�yRHXc�i�u����
�'�T�
#��!Yo(�Z"�2h]v���'>N�#��
#@�Q�L���H�yB����� 8#�?5�L�@R���5}h���.�6>��$��	Df�ħ�y� bK>�ç	�N���ԹF \�9��ċJ�I��Tm�K�M��ӧn���'�$>-����/�z��x&��ɣE��d8ʧ)�Cq+�6\詐� J
QL��mx?iӥފ�)�S�+e����^@��L�4�2�B̐;< ��|�V�ɔb���S�O��$��eAp@\8�쌚uz��!�R?�Y~J|&��S��U��;S>����E�T�	���,/��$>��}�Dœ8x�Yф+W�1D~���)�JU�#Oq?Sħ���� �5##�/$���Q��ȹ(���ieqO��S�O��Sx�0j����u�z�ȥ�߮Q(lc������R��g}"�I�(����FN�$)�0����������<ISVep�{��)p�6��FK0%@x%b$M�(��D�(k�6[�{��)�s���A[�à���
��D3�����	�8�=�)
6d�>+�E�`�HZ��B�GC�9�GxJ|��d�%��A��l,@�#�/R�'�Z�����ĮHhpy�D�Q�Gn\�	�6/ �ɦ�X#<E��-�/E�Q��!5:��k�,�M�� B��c�~��~"��$�
�"�q!� �*4QV�8"��9d��d�'i��rad
�s�a��E�/���g$�-��� ��-���@j���Ä'��S�O��篈3*%�� ��D� �4@3�'��<�B⎍"�J�O?���''��I���YI}��t�o}0�y��݄M������Oa�j��u*�ȺA���S�� �bȊ\��Q���,����BT���SG��[!,Т�>zp/�;S-x�y�G�<��D�{�ޝb�S>R��!U�<|c�/V1F0����VPQ q�i���"�(�Q���"2�O�<8� �z7�x�C�A�}1�'P�Գ���c��<1e�@(�!0 �
�^�M���A�<q�˞@5 ��T�p.����}�<YA��?���'��SDUz�<a�%[chE�P������~�<ф/�C�F-���]�Lk��{�<�Q�-d�8ԢD��v+p�t�b�<"`�+1����Y�n8"8
B�Ca�<ᕠ��
� �%j�>�nA���_�<�G
S,gl�QWkɼ���)2Ob�<A���
�hHu�[<6�������E�<9�#N����c�73� �t%X�<�d+�=g�>�
�J�S8)���Z�<��$�F@i`B9���j�m�<�U5l�z���W�^��A�G`�<��4R��@��딭k�}k�b�[�<����O��L�D�F*�,�P�ˈ[�<q���4��Ѣ.]2p8KF�RX�<�V��m�F��Q�G9?&PHq樀j�<ᡧ�)�R�h�c����5�}�<�Go|�Z<�@CZ��m�Q���y�jԎF!�hq U�� �A�JI��y�[����v�6#�M�R���y`�A�8)�r�*8S�a�y��ٴ]�<@j��2y��@���y�L��lyҳ�5vG:TB"��y�b��.	���._�h��$٢Đ�y�Ց;��|��d�3-t����y�!R���u��>,��Q���yb�^;b�%���jF��$�C3�y�bQ��j9��s�i���y��h���A$)�@�r(Z#L<�y2Cs8��X2�,ԣ	ێ�y�mBgd�%�T�
�ts�pr��y!��,R@YA�'m�������yR͉�e� ӗ�ƅ;)Te�z�<�&ҙ=+�4����\𧍒U�<�`Ѭ'.����"Mpd@`�LGU�<���Pܚ S0M�
jBu��i�T�<9��ͺA���zW�2Cn�VC\P�<�&O)�|���۫!~���R�K�<��F�kx|pE��	�PkD" K�<i���*��jGI�sG��
�
|�<��E�6dK���F��Բ��w�<9q�b.�$p�Iİv�~lb�N[p�<���
�`Q��(%nٯT����S�<!@ax��1
�W�K�Ҩ���_F�<�@�#T}zT��c*y�b��§@y�<� �Ј�a��) � ٶɆ�6k�EG"O�]�L���(�R���(,H1�"OL�b�ѫO ���v�P���"OY[7ĂL݈�{7�Q �6�:W"ORmR�$&-pu{�C]���[e"OB�)�J͘98�C��(9�s@"O����>��3��<�t)kS"O���sf��vh��f>�[8�"Ot���յ>7^�[u�`�� �"OfI��#�d0�C�HܜR�ꈪ�"O�E���4*�D�Sh�	}�\@#"O���N4%�.�1�i^���`C"O�
�)QU�|���²��(YB"O2�[��Ν5�r}�
�$�z�A�"Od�3j�;}>�ӒB�a
܌S6"OF�	�IƜWVT��AڠR���r"O�i#��݆i0bV�[/]&����"OF=q�d�<�|���T-4��Z�"O�Ԉ��E�c�v�BBO� \B�Ib"OVx����v��P��:�\�'"O|�KtbC<}
�`�I�Z�|iڑ"O�f)Y�r54�� LӖz�-"O
�*�`N�x�(�#�ɓf���"OHI ģ� N�"�h�+�@��'"O���#�:zr8P'0-���"O&�YGL>OB�������T$�W"O �M&aS������"O��#s�^B΍)cH�D�<�SS"O�h�M�5Dl�b�Ԗ@�z,�"O&-�����!v{�F�+ls� ��"OʹCR��$i��I�E�@�.��"O!
p$jP��s�B=�e��y"��}��E����3\�QQ���y��9C�x�#�����A2L�>�y�M,Wp��v=)�n4�aď��y�^8r	q88�� ͙��y��T"YM��в�W<5U���@�y�O��w���`^!'��q���yB���%�B0jf.�	2%҇C[�y�mg�D�S�/��~��M��G!�y2*Ƙ[��h�@ѵo	� ����yN�2f9̡��C8f��=S���
�y"A�"X�5i�kϳV����!�y�g�[�,�JAO�<�|xF�=�y2�K�q3޼�ߌ�y�'ɘ�yG�q��m�D	�{ �a����yB�EZ~*0�.9^, �(��@��y�܂1ƌ:��S�.d"��L��yr�Øb�0�k7��8JP
��e>�y�eݷ�$����I��I���y��H.}F�QC�N����kS�X��y��v�nHK����LN�\�R]��yr�I�,�ʌ��������a��W��y��AQZƍ�a�Ǿ��������y��G����D8�,qa4 �5�yR�@%\���Ǧ�?�lX	q +�y�I��|=��lɈz<�;����y�!ζogH�-@�k��uYW��y2/N�	�pz7Aձj<�yc��y��'z\�Y�Ҟ^����,�y�a�p6 ��S`Ϸ_%��b�*���y⢙2�J�� �ƫR^�I��AS��yrʛ�M�L��ҋ�Tt��l�>�y�A�`�%z�� �	$rܑ��� ̸���
+I���ؠ
d��&"O6�hq&�z�i�p T�^�p�c"OF��CV�Y�N���W�vB��[T"O6�y#�F�cs�p��l��u�"O��Dȉ�$u�y3-L�{��i��"O���L�*�j}8�@�bm���6"O���EA�`Ų�P�Kmj�X�"O�L�uJ�&�����+6[6�*s"O�2�*ܭSOƥ��H�) m@��S"O*hZ���6V*M���T�p[f��"O�[<>�0��TG������"O�]�Ć�"_���D�(�)�"O�-�FO5V)���`>�A�`"OJ�C2���������c7j$cb"Ov]!��!��B&OՓ(<Q`�"Ol�`p�,-?�ͻ�.� 쪶"O"��!�l��43o��!�"OJ��&�F.N~н�e� ������"O=�BY
����l��u�ԓa"O�e��T4R7��	F2K����V"OxTh@$W�!u��E�I+w�e��"O�	��;a�x��� I��(1"O���f���3��e�g��;�-��"O�!���0d��U���݅%��Hc�"O~��d���1Q�`�׭N�!��"O�Z���dN���G*%���g"OZ��`!�H\0i(�d�r���'"O~��㓌`��P��j1k�2D��"Oȕ{v�E�Cl�%j�;6հ�j"O�����r~��+ )ݣm�p]�"Oj���A�,/`�1�����h"On�XDmD�|0а�F -���"OT���^�>A1у�͢8𖼢T"O��A¡�M�x�BH���e""O
 �kǲG�x�i#&Ϭ��� �"O�Y�@O�D@�-is��1a�Z��"O�M(sLB�5Ւ�#�d����1"O0
ը*�p��dˍk�};�"OB�I$�
c�έ�Хϼ�T�Y�"O�ؒ�
�b�@�ŃC''���b"O0��b˰�	�F�8C���"O>�X��D�W ��j�<c8e�"O�AaCW6&�Imm��<��Ӓ"O���%�)��Ԙ%IV�=$���u"Oh6ϖ�+�ԉ��b�$:(����"O��*5j;V���A�͝��c"O��� '��\)���R(��"Oj�:�eO� ���R����a�,�k�"O�u������#'I"�ʑH�"Ol�@��Y.�0+cރj���!"OV�eMݾf����D�c�Jx�F"OX�aǜ�:���!A0[/T�±"O�X���1/+츻 �#Lʵ;d"O�8���ۺsj�h��i��)Rܙѐ"O��J?D�T9§��I��d"O8؂B*B2S��%
�I�G^q��*OZU��� }~$\Qa�5.��#�'�&��X��%�Ӯ��n��Z�'��M����l�,!3��/TE�'N:u�sƨW��]�� H�x)R�')��a�./�T�;�C�8����'�L�%���B��%���&}G�l��'h���H����Q:�,v�=��'4�Xi�ÅZ#r�
�*�9uT�K��� �g�R+Ɉ�"dM#/�����"O�h��������C��y�8ႇ"O�ո�	φ���zc���MP"O
�Cb�� <e�t��!��m(�"O8���`�!/2>0k�M�.���`�"O��5��7)� &�
#O����"OΨ��'y�ƨ "�J+$�.5�1"O��;%O�0R`Js�V�#.�@�"O���F˼#�:�K�
z�Ȭ�""OJ@v�@��
baZ#x�jy�B"O�LK����@�v9ɱ��z�A)G"O~�KR.K\,��[�D�}1�"O�
�R?dK�m���ٸC�uj�"O��r�B�O(dأB��5^�k6"O�-K�/D�G������GC��s"On��'"\*"����f�RRv��P"O����Uazp9dHϲxކ�je"O�Ū�J'�L�ʶ�Y��4�7"O �9A!��{k�U�q��Z����"O��!K���
E%�:w� �W"O����.��-]:z�ʴh�"O(��g   ��   B  *  �  �  �+  "7  �B  $N  �W  a  �l  �t  T{  ��  �  /�  p�  ݚ  /�  o�  ��  �  4�  x�  ��  ��  C�  ��  ��  R�  B�  ��   �   �" �( / =5  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�Ik������@�d��M3��L�R�f岆�1D��ȃ��m/,�Ju(H	|�,qZBɰ<�
�IL ����|��0!)�e�ư��6ڎA�7i�=z$}���6 �X��a�����.C�#�(`̔44��PEzr�~�ūژX'00�N��䕋�%{�<�@��`=�� $@	�D�j6΅Φ�E{���i`�!3@�)�*��u�W-RL݀	�'�\$[����
���G'"l�O$��$ڃZ��㓂S[)ʍ���C
�!��Rj� �S�MH��B�t�!��e�X���D;D�R�qV�D>S�!��Mr��U����d����P.A�!��'	B����]�-e�KCd!�dG*}����2�����	��1F!�d�8[㰩�Òg�X��'W�j!�D�sO�M�� A'g=>�;v�X#:�!�ď9�i�M ?���� �=
�1O��'w6"~�gJ��H�5;�-��@!g�]�<yS�۽&ę�ċ7*jph���?�a����FE	�6�M`�ԛ~�;�U�3�	D�B��A��'D�U�ȓ&��ʑ$T�[� �)�I/9H���
�M��''�'���g�[J\P�D��s�L�g��8���'a��O��>A)5�'�l�Iᐭ�*�3S�/��0�դ�H�!�D�4I��� �B��t�j���m�!���J���#t�T���[�ni!�䃻5�|��R�&h�2��`��/a�� oR����>	��ɶC ������A��,��^|�<� � � 	I&/�~�#G�I'1f�E@�"O�aud��D̼Q�@�cf6y�s��dEy����O�PPEJC5A �(L�7�Ya�i���ϸ�P�d�1{�2���H�PV�q�����~�1�/��0��M.i{Τ���O(<9�4
1r=�'�@(\�8HCQ�1t}���0�|"$,\O@�	ť49��+�k�P�F����'��O����k���:�����y�"O��r��)?�\�6i�wς��ўx2�)�ӑ9��"�^�<yIă��7�!�,ɣ�ڱ�(�P�+4R��q�8D���D_�s��g_�u�C�� !���k��4C��-�Q#d�I )j!�䜟(=�srʉ8X���{�DՒ!h!�Vw-�!!GU9��,Ze :#f!���xΊ��$�A}�XL���]M!�D�
�6�D��AL�K����mQ!�]�76��R2$%h���7*!��ˮy����d��Y�\�)�@׵��y��I�C�>��$ٯ<6�ph2�� �.B��,D�r�����̐��h(yU"O
t�c�;'수�R��\@�X�"O�,:7�
?���A EP��q��$~Ӗ|��I?I֌�$C��~?��m);�PB�ɛ`����#��)C�Ё:Q�5~4��D+ғ74
�SW�� �NŁ�ǀ)ur����ɦ	�'��	�|�qq�#J�j/�KbϾp�C��:^e|�b���4o��`JgAN�La}��\~�I.p�<) wb�!�`���l
"�yR�M�S����'���A
"�O���B��	�<),O@�O��AD�[�ԢQBF��>x��'��	�M#���MEܤ��dE5G�]��COy��'��v��~e$zD>�ҥ��{B�p����*�O�6�9�<�?NT:�˧�\��!J�$��D�x�Ɠ<:��.ǥ��Y9��q�D��O�6m�>���4���k��v�(��I��
�8D��I�+2jD,��!h˺_8��G%#��O|H�y�K�>��O�y@E�C��ڡ�Z�nP∢T"Op58�h�$�\��G��,x�ܤ�P����I�FR��׫��0�ɱl_�jN$C����-��H�Ԇǘ[�C�	� s�t�!�X	�2��}.�O�=�~��MKC��c�+R����I�ܟ�'3���$@?b�㢀�'�`��t(�6\���0=��'�JD� ��<T�e�g����)��xҬ�)|���`���Un��b��B��y�����ȓ��H�I%��HGր�yB�
�i��	�B&p(̌��G��yrgU+.@���H�2p���j�e���y��_.4�p��ij�j�z����y"Dؗ�"�Q�-�[��e����/�yBG�,(;�P����i+r/H�y⎞;#�����
!l�!���� �S�OI�é�%w$h�k��BѠ
��hO�U��/��k��� ��Kc'���$"Ot�2U%ϙ.V� c�#�&�R"O��{e��s5rp���3k���"O�q�&@�9
H���Uhc��o�@�Xb�C˕v�����>�N����2D�<��sV2%�ʏOHfL��Փ�hO?����w��pz֌��?�8�;d@	"H!�dM� Qa��7}么 K�A�!�đ%p�v�`�b�qo�ա�% ��|2�xB�D,k��K�&��0��".��y
� �yRԍ��tL|2f��"y"OR c�@=�n���O�K���X "O8�;c/T��5�vgȝ`za��'�qO���N8Y���z�蜌k|jax"O0B��8`I��'&֤c�>��]��S�I��#��Jx�JGكj]����'��4���΅�{�����ahX�Fy��'���ke���, ���10m��ˍ�d!�'|�*1��׹`jF|z�g�/1�Nd�ȓ�*�k֏�.@����+_.>�l����?�}��i^�|4a����/4n�`��"��C䉭r�^�8bě�H�f��qS�E�Oh����I��;��i���D�8�� ��U��!��9D���`񬇇e�<q9K���!���f��U˜4P��yB���;�ў@D�	˴pS~h8M�*��ti%K�j�!�B�K1��1d�Avnu0��)m��y�	6&��p&�=�Ihb�Ɠs�XC�I4��R�-Ӣ=�@��JC�Ib+���D�5S5M�4q(�����>�D M+r�������DkC�Gq�<`��fc�ݫR䋨't^�uj�a�'��q�O,�P�%&�	�a�4gI�z��
�'}q�jO�$�lXy��	+E�葳�'	ў"~"aMƮ�dt����r� <Р̔p�<�vA+��)bQ�S�{>��V!�o�<Y7+�P���Vd_,pK���e�Jl�<��	�4�n�
��(<�� ���WM�<wc�<����n�e�����JL̓6��2�4�aDJmr�5acEZ�� "O��0l̦8�r̨AǙ=;K�I���_x�L��#��!RQj����{��x�Bf<D���gdY"Ġ�F%-D�p�s-D��C&��9 "��9 /�����e�>D�1�j�1B)�0��ӬE:�iBF>D��24�G�(PP9��G�-n�p�'D�� �V<�Ts3ZA<A�&�*D��@���qԈ�SIڨ& ��gF%D���% �~�r���H�>`��x��*$D�)��O>RuD���J�X��� H,D���T�B�f5b��"�PMZl��a7D������@U������Wa����4D����Ƒ�
Ä}�I �t�ڭ;t�'D��@DK��cb�ɀ"C�Fj'�&D�� "J�!�ĩ�Q��=d=h�K*D���l�z(��{D\:M>5Bu�&D����C̾D{
[�1O&�3��/D�`�AK%.&�
��W�o��	�B`-D��S�/� �����e�xP����*D��C�j�!Q��(��S�t�΀�#D��1ŉêk�Z��A���bԺ��d.D�\#�'�,]�4Y��Ē
��0I�&D�H�g�;����@��!5^��Ff:D�pXp�$��"pNv&��d$:D���F'�+�Υ[քܪM�����*D�li�	�O4Q���O�\�Ƞ�4D���c���K) �W�y���b��&D����S.#Z�}㧈J����օ&D�آ�;W!�TEhG�z�����J%D� �A�Ӗh3"��vCG�d1��Ѐ�?D���$�że�)2,D�S�v8�w�(D�PX�B��5��@sԢ̈́,�8�;pA%D��i2CM�q28�9D��5�F�c�E/D����,px�8���$#"E��-D�� n��ץA�L�~A�Y4_�^i��"O@\�ץBi�0qr�����bT"O�����4!a*uۓ M2�#A"O��CA^�Cs���M�9HJ=RQ"O4(����p�00����4�8��1�'�"�'���'u��'���'�R�'��Kǟ�_�^�b#���Ta��'"�'���'�'���'�R�':����!a�b����C[z9i�'k�'y��'j�'��';B�'Y�e��ƆGIP�ɢx�0YV�'���'���'R�'��'3��}榰��A5b�~E�ѕ�h��I؟���՟��	��T�I՟D���$�	�6�l;D*
4?xJ�������	�� �I�P�	Ɵ�������	П���(}j������ �^쨔�
O,%�I៰��ǟ��I���	Ɵ��	ٟ������ �:&x��hS\�8���ʟ��������h�	��p�Iʟ�I�BF�iJ�!��y�0E�SLH+P@��� ��ٟ����������Iݟ��I�[��(�G\�6��I��L% ����ȟ����t��ӟ��	؟@�	ٟ��I	o	�g�(=�f8H�O�%�8��I�|�I͟�I���	���Iӟ��ɬT�"���_�]� I���h����ޟp�I���П���՟�Iӟ<�I�OJJC�.��h�@3b*	J�d�I�	����ǟ��	��9�4�?���=~��S�K��/Ɩ)�2̘�:ڢ	�W���py���OxdnZ0f\�9#O (�¬2 �K�f3>�Ç5?1��il�O�9Ob�DC�v��!
���'L�T���$3����O��Y�H{�j����)�0�O�ՈdMO R���s����mQ�y��'���u�OU��R3����>H���I	��v!`�Ѣ��*�S7�M�;JǄ5C���x�$	� ��q�"d���?!�'�)�Ӆ"nHl��<�p�F�|5
��$iB�U�C�<��'��	�hO�)�O:P����it�]�E�u�|){T?O�ʓ��
p�v�ڎ��',�9��d^�9��R���UfX����dIx}��'y�=O��Dz�툗*&�X�#V0R]�'r�8E�6�j��t�C���j��'��A�M��afG82p��C�Y��'q��9O2lC�A<Waq�!��d���F;O��n�/N%`�����4��`��	��H�!G ^z���9O��$�OX���;&�F6�/?�O���	��3�2���c̽/@���_�8}252K>�+O1�1OT ��K2Iu���dCy��4�S��P�۴q�����?����O�صbD<b�X�r*�*�����.�>9���?�L>�|Ra̜�a,��{�'Q\���&�,�X 	�⋆��d� r�lC�'��'L��'V��ywȇp<h��D^fF����|��̟ �i>і'p�63'8�$��{�l$���\�L$Q�Ì�C�����?ёX��	ϟ,�I�
6�h��M]5j��u��i[2N�-�%���A�'�8��f���?E�}���}i�Pʶ �j�����-�V�B���?I���?���?)����ODH��V�P�Q�!�1Ɛq�Dja�'q�')�7-Ҳs(�	�O�-nZH�I�[2ez�+
 H��1��"Z�yt�'�0�I����h��k'?�wK�#;��ۄ���A���E��w*�T ���O
�L>+O1��;�J��� ����j�6l�$��4.����?q����O�v�Qj���Z��m;d�s��	�����O:��<��?�X��O�B�t́��0wf5R�ыY��إb�xht)���C�K?N>���f��5� $�+C�D�k�M���?���?����?�|-OnymZj�je+!��;9�jrj�	jz����V����	%�M+����>I��q6胢�M�#.�u@'$�ԉ*O2���&�	f�IMZj5aq�O8�'�z��3
ݹU����IX����'��IܟP��⟈�������b�4���H��چa��$��+��7�Z�o�t�D�Ob������	�OB�DU�� Ǽ�U��]���jF����IҟX%���۟��I?� 9�`��(��\�!�2e06B��\�lL�i�<b+�c&�͆D�ICyʟ��L��n��h@��O'���[��'@
6m��s���d�O���J�B���AI� �PM�E��\��O��D�O
�O∐wK�+�����2E�P�1���A�ѡ�^-#�@N��b ܟ+3f��t%M�"�Эi_6Q�c������	�������|'?����Bt���~G��Pu����CЧ��p�n���M�rcZ��?���֗|B��ywMU8N ΄y�Ï�#�+���y�'�R�'�Đ9 lU8�y��'"��+��]�?���b�GB���C
Q�tۂ(:ÍB�f�'���ٟ���㟐����h�	E��8�DP7uU��PʾNa|�'�H7M��U"����OR����>�I�O��C�UĊՊ�A��̰�DT�O��9�'�2�'�ɧ���'����wp�Qd���^�����L��nH+b)�����o9Zو�'��'��	�Zl�Sg���b���O{	x��	�����П��i>�'b7��=38��D�,�P�3cK��=��)��9v)���9�?)�_�����)m�j ɐX��I��kM��F���@(���3=���%C�4RI~�{�? Ua�d��x�a�t�ŋAh@��?O����Op��O(�D�O��?��O�m�p�ӢY: ��س��ʟ��	ğ�r�4!��'�?�ѳi��'��dq�G7)�c���&������|��'7�O��%�b�?���ߓ.�y�0�ޛ��p�blՏq2V��@݇�?�7M/���<�'�?����?IfIЅb���c	I.n���gcN��?!���ަ�BO�����	��ȗO�V�;;��`�Z��j� 6?�P�@�Iퟬ'��1�^Ih�ǟ~ИՈr!]Z(�	C��̱��s~�O=h)�	�gP�'**d���P̕r�mA��	�'Ir�'�����TW>��'h�6mx�h0�KH<pSmf�Yu���O����!&�����d�O���ܨ;Ry	�H�3��{@�O���щ
G�:�1O^�$ܨ;Fq!�'1��Jy�mѐc���PD@�%b�ϓ����O����O:���Of�$�|��OO1z��I�쐌F������j���J�9���ğx&?u�I��M�;mb4�b���(ą�o�� ������O��\R�h��yB돤i���
#L2B���y����(n�%��%#}�'k�	ߟd�IR
����L4b0�푀'IL����� ��՟��'��7�R�/�����OB� �73⩳��7!�q$�'#⟰��O"���O�O�ZN� N��뤣��vW6,����p�wLǞ~,FxQ�ADF�+BAԟ,��'�o���{��J��(!֌ D��h7j�

@� C�$T��@IΟ���4P�ظ���?� �it�O�nI�zr��e�7C4��ᡉ�	��$�O����O
��2J���i݁��?���g��ZE�'�ۓx�@#�T�l7�'{�͟0�I՟x�I՟L�I�!���"$Y�I	���e(
�X^�a�'G�7�S�sU��D�O���!�9O�|jw0+bn��Q��5����l�t}r�'}��|���oV��J��5Dl�`���@����t������)D�z���CS�Op�9�vu#ƍ+\��8�b�0�a��?a���?)��|�.O��mZ4 w����*x�T�5ș�!��1�����fxȠ�I�M���!�>a���?�;Z"�ي�G��N]r�s��p��!��53y$��'�F�(
D�?aRP��d�������p�����;�+� �yR�'b�'���'$"�)B��zѱ�
Gg����% M� �$��Of�D��
u�v>��I�ML>9��v�x)x�
N9#r�cB����?!���?�͘��|̓�?1�n��Dt��D#r�|���ϳ7�Bx��*���'�P����'|b�'�$ٲ�㜽w�=��W;\��H���'RV��;شS���B��?����Jb2be���&	�;�k��c������d�O��d6��?�2���)>����cF�u�(PO�/���BB�G�<f�锧��+	t?�K>)խ�M�&=��a݂'�"X��	.�?	��?���?�'�?�������䦑Z����5���0��� 뎘+q)U'~$!����ش�?�)O��R@}�'�����4��I2��eI!H��'q��ME�����'[r�� ��]�
��d�c�p�"�+_.q��E*�
A�2W�$�<����?��?	��?�(�@�;+A�mw��(�Umw�}S�C�РW��OV�d�OR��T�����]Fj\�r3��$$�$�꓊�/(d��	J�Ş|l��!��<�%e�^F��Ps"d]
��E
�<�e$Z�1%���8�?�-O���?)�:�����EQ[��|x����yx��?i���?�)O�TlZ1F&6H��ϟ��	�c�0��FY�"�T3���0Na�\�?q]���I��t'�X(��~El(�TC��Ԁ5Sv�p���N��Q-۽e���Z�#�O.����W�|a�d@�##�h���LoJ q��?9��?���h�P���!���0V�ęd�\�f�ǣ v��ۦ��k������Mӈ�w9�"��ƶY<��E(2'ni��'���'�R�N/oS���O��Dc���zD���w��8���.���酄+.����4̏{8V8�1�W�T\��ҨL:Gפ��F�>� e��!:����ʮ3r�Q@�˳B48�)� R&3�P��@?p`�J�����Ǵ�����nlh	�1Cը/�>�s�#Z�#���Y��(f� pW���j��a��b���r�}) H����,��XA�.�;[��0ց��R�]�S+>'c8��ʍ?,9�fZqɪ�q݌V"xl�� 9s����-$;�}d��4X�yrd_e��.��m�ѮW�h��F^6����cfT+ �����)I�_m\q����?!��?��'��$H%	�9��j��|
���'��$a���m�����-:'(�?�~�/��\8!/Ƞ@�r�ަ�łğ������I�?Ŕ'�b�'��<
��8ED��6l�Zm�,i�<��� �)§�?� �CL��h�^�z��ORCZ� �4�?I��?�7�����O����O^�	�+V����X�S��ňЈx=xb���TE�O�I������Xud;p�&�*&O��(��`���ܐ�MK��\=J*O����OZ�$-��Ɗ�A��^��P������<�@fR�H����򟨕'��'��V��C�-\={\�Qg _�Kt��X5��ٕ'���'Tb�|��'U�e�Db�X񡄦7+�lS���.Y�B�q�y��'��'��0�n��Yd�q!�V�ZQ!�L>D�Yl�͟��	˟�'���I˟4�D��d�c�y��(8T&U�Sa�y9�����D�O��$�O2��r��,�:�$��z��)�g㋰ �i:Ό�S>�oZҟ�%�x�	ҟp`f�&�)� f�F�f��}z��F;0��Ek �i���'��I�ro�	�O�R�'����F�I��mJ��T�C�0$�Ov��ObP(�k�Ob�O���]�b�����	>N<T�vh3K�p7M�<��!Y��?)��?i��b,Ok��d��u���ݗ:��Y'�+:����'B��7��O��$�r�"[k�b� H5Q��񩄹i�T"c�|�0���O(���\��'��ɷ�d@l�!.�ؠS�J�(}mFAa�4w<8(�2�	�O��a���-I}�T�Uv�����/[ܦ��	П��	8>G��'E��'a��Or-	D�L+�~,y�c�M������R~�O��d�O�=5�ց��O�#�X��`��P�bm����Ӷ��cyB�'��'�ɧ5VM#А\P/�$�Ɉ�������s���Ox��O��d�<���� h�m��!�	^\܊`��:9�\+O>���O��D(���O��d�g�#�Ǯ?N�����{;�*�H1���O����OzʓD.�� :����"+Ү!�
��1�N)*��  �Y��IޟX�Ixyb�'x�2�2G<1#�4����w�:	i��ՙ)���?����?.O��â.�g�S�'�`�ٳ�Vϸ)�%�+Pi4�`�4�?YH>!)O��O�O:Ʃ���[�J�h�2ŃܨAT�pr�4�?�����$-�m&>��I�?ט&}۬���F�
cd�q�#�i�7M�<)���?����?J~���!(/���B��a~.-q7.���1�'@4�ڳi���O���OÖ�v�J�!媜�S� ћ!
�ͦxo韐�ɟ ���	����O$�)�|n�.8޲���E
���c(Рb&:�48�����i�"�'���O�O�[�W���K������;���hAh�n-
(�����4�I�D��u��'��_��20!���cVv=��Jŝ;�>7��Ox�D�O�P� g�i>��Ɵ�ˀ
�h,A �H�0)<�i2'�M����?	�������Y?���I�ȁvB\A8!H�j�$j$�8��	�M��r��Y�s�x�O���'�I\EX�f`��Z�ig�n��ٴ�?��-���?�*O����O��ī<�3��� g�r��V� 1�KQ�S�J\JE�x��'���'/�	����	?]^ɳ�G��t�6Q�FnD�Lb��.��l�'���'��IşY��Vx�Z��\�r[�V�2qFݫ)��6M�O~��4���	�6ՠ4�)vӘ:@��z�����ʘ	޼�3�xB�'#���d(���]���'H%��@8h�]:�hV����R�iӢ�P�	ԟ�##fS&� Ol�#��4qp|��O�l��Pói��U�d��!'���O���'*�\c������R��2G�H�����M<1��?�����m�<�O0�l���F�.��x�F�N	^�p�O��DF)|pL�$�O���:)O��F��T+�m�/ƪ%�MM�cn���'�b�["j=@T��y����.m*��P�Q�`t�I��N:�M�b' ��?y��?)���"/O��.zV���L4[6�k*AMT��ݴ1��:t�Y�S�O��9�e���j=��H�NBq�'�w���d�O��48��S��>a&ʒ&�j�X��q�����]��:����'����Ezҥ�j<[NP�6���V�'ΰ]�w[������,�È���L}��$�y�83�
���N6��'�B�'��\�,��DL[F�A5�ģN��|���jB��L<����?����D�O����,c��ԡ:R:�˳	�?��1Kw��O˓�?����?Q,O������|R'm�-R�e����.I�e@�l}R�'���'��	�x��t�����=[�:(�v���d�
8[��2-[D��L<���?a+O�� �r�S�m��H �(Y+(m"՘���!�(P�۴�?y����O���хM�2�d7�Tj�%pnH�!��*P����W>�M����?Q-O�(f�\R�ɟ��s�!RS���ȑx��]�I5JP |��ʓ�?��g#uI����'���vZ����SWh�뢣�y<�mKy��B�n6�HY�4�'��d�!?y��ܽ1<x#w��-"|�y��$�צ��I�)'�F��P�J|b����iR8��g� 3nD+���c��mP۴KA�tJQ�i��'��O����'���'Z�iVd�wza91�]�"�x	��Jl�I��O$�ĵ<�'���?9�fG,��i����:�,��s(:S�V�'\��'�x����>�*Ol�䳟�He�r3�A���V�oy���#uӀ�O|PT4O������������W�Emv�xa
�0&��a"G݄�M��M��U��T�l�'��R�h�i�=J &Si��(���K����'�>!��J�<)�Ӳڴ�?1��?!/OܕX�MC���L�t'ԋ
�����VE����'����ė'�R�'��T75���@�j9U�� s`�jY�X��y��'��'���2Do�Œ�O�(an�b��Si���L��4���Ofʓ�?y��?aBJ�<�$l�>���H�`��:��ȽQ���'���'"�'~RfM���6��OT�Ď6 C��r2oD�?)�Td�<B
HTl�����I�'Ց����'%�d�#+���3�n	$H����R[���'��'C��E�7��O2�d�O���ȡY�((���_��> ����W?�mZş�'~��(��D�'�i>7�մ�2�!�Ύ�Q�B�B��59��&�'�R(��[YV6��Or���O��)��N���5i=���"�E�Mn����*||�'-�V6�'k�i>9��� `4�ӏ٣~_ĔC�nq�m��i���RĂk�:�D�O:��䟨���O8���O�����;����5��43����A�����i�֟��'���'���?���&f~�R���/+�H(��_=Mכ��'B��'	�y�'�z�>���O���O����ta���8o@��P-PT��	��in�]���Fm��'�?���?i�b�&h
����%6�*��tE,X��'��řD	�>�-O^��<����v�>[��	B2���.(�1��̀{}�R�y��'��'�"W>�	� �(�p�K�:��Y�1BUod|��G����ī<������O�$�O:l��	Rlꐘ�J�W�h�12ā�����O����Oz���O��<�N1W?�$����-8� �r �.�L��i��IΟ<�'���'8R�I��y�o1b���蕈��JT����N�a����?1��?y,O�����u�t�'��=x���d��a7����[��Xڴ�?,OB���O��dę,�1��v��0�X���؏*��gV��M���?�)O� �B�X�d�'(��O
��8��)$�Bc��% q�Q	Ӧ�>����?�� B��͓��9O���r�-i4�B�^�N4�TC��7m�<	���%xћV�'{"�'���@�>��8���g��.mY�qG�9{�|�o���ɱ]z��	��'�q��NMb�؜B� K��`�c�iԶ,�`{Ӻ���O����a�'-�IpE�U�7O�j!���w")-���ڴLSTLΓ�?1-O,�?��I�z"$\	!��^;�؉G.�{F��ڴ�?Y���?����/A��Hy��'L�$[�4A�Y�A��ݦt�t&@�'Ǜ��'����(�)r���?��4AX��&��(��@D�V4"#k
�Y�I�1����O���?+O�����L��˂@u.�hfQ�#�@��X��;!�`��IƟl���d��y�fF)SčY�L��H�r�%E��*�>�(OT��<����?Y��k��`c�R�L2�"i(
�A�h��<�,O��D�O���8�Bs��|�GM�m�ޕ� �ۡ3Z�ㆋ��	�'��[���������?a���2v��u H��H��3�	tP.x��O"���On��<!C�_kv������M�1����kކh4��Z&��M�����d�O����OA*�<OD���O��ӨW�G+<mxAe
�kki{�/���I�H�I⟼ku Q�M����?���j���3T�v �ħ���R�R�y����'d�����+�jy2Q��s�|�p��G0C<�����00ߢ�e�iOr�'��(V�{� ���O��z�)�Ob��vB�ib�a�U�7�����D�v}�'�f}A��'b2�'��r��B8t�&y�B�Fi�s��6ԛ�ᏼF^6��O����Ob����|���O��1;�#j_�,9	��
�~@oں|�:����P����I?���Ot���̖�H<���2���p����������I<A��Y�ݴ�?!���?���?����)h��A���4���8h�en���<�'.������O�ĺ?9��
\�EZݩp���B�gq�@�$-6b�����`�ɇ������RGE�E�����T
ѓ��>���`̓�?a���?����?��e���9Kҫ�C����E��Uf�tH��iH�'S��'����d�O�P���R`��/'Cv82�`�Q� ��'�������L�'rX�	�i>i�!V^��e1��D2%�P�᫥>����?�I>���?�aP��?�K'm��`��)@��I�L-&������	�l�'�N���!�i�%p�zh�JZ>w�L����{u��lן�'��']����yR�>�셏u=ݸ���=K`��L�ަ����ؔ'C�4#v�'�i�O���$8x͛���'5Db]aƀD;{��&���Iɟ$S��n�`&���f��V�Ϧ?;pl��L��g���n�Ly��f��6�Ik���']�$�(?y�'vt8	���R�-w>d��Z�!�I��
��a�L'�b?)�%�0�EڃB��,�T\(�dtӶ�t�B�A�	��$���?�sL<q�]�X�v���W����F�jx���i8����'�ɧ����=���K#jJ	���ЕN��. l��H�I���*�g��ē�?���~�ͱ`����]�J�Ѐ�x)n�q�ɵy�=RL|����?Q�O8n����Sb��!��kRhܴ�?aD� �5�'B��'ɧ5&kG�X�kV�԰�dJFJ����;��İ<����?L~
�"���"��t��!x�aPQf �-;w�$�O�OV��O�����?k��� $��Ĉ��@8R�1O����O����<���w��)�/��hs�ՙw���F�e߉'�2�|��'��S��D�Bjt@�Cݴ��,s�jԲue��۟������',��.Z�O�.��ɜ	6�*!��� #�FyRp)p����5���O��dS�'N��8}��P)�D2-�aH�4����M���?y+O��s4�IC�S��S-P�1���E[b}��(9�K<����?�ō��<IJ>y�OuL1����M�l2e'�v�ܠ�4��$[�|&�oZ��)�O��i{~o�$�<Sf�ӘN`�&�
��M���?Y����'�b?��$���AF���$Ҵ,���h��v��:f��Ѧm�	��l�	�?�)J<�����a����*q�ߡ��%9B(���s�@����'�"|�����2�C*� T�2Ip�吠�i��'�b�%�2O
���O���:(^,�0�ġ��c$
�#�7-%�dGr=�?I����t�g�? �$��Ы4�V� �G����E��i��.��O����O�Ok����1a�$��UÄ�(!'S&#�I>f9ء&���	���	Iy��+9���ұIL)#�,���G�EAbջcg:�$�O �=	�'��8�M�p�ԡʹ��d/5�b���<)��?�������MHb�ΧA����jڦ`_�Uw�D�'�"��Dy"�'�N���g�8l��T�eh]4-2h�ہ`�>����?�����dXg�ܠ'>�Y�D�?_�H0�%����w�ߖ\�x6�7��?��f�>�?)L?0'�Hƴ����-�0�Ok�����Ox���O�<�2b�|����?���01"�ItW�!GN��#/�n�ZP�x��'��Z�0vP�y���5�Hȥ.���֦1�5���iR��'�J��dOf����O�����|���OkL՜���p���Z�y5�_���')�!ڲ�4�\�'�j)��N2c�"�A��; M�ٴ;M�����?*OF���O���<�eO�D��� UP�iQ��
5����0" ���y��i�O 9���/�����R�6�VMH�c��5�Ivy����q�Iwy��'a�dڴ:{�z����m"�(�9:�X��<���E{�O�'�Bg��9D*�'4j�,ce��0��6M�O����F�Q}��~���?9H�3�N<9q�d3Vj�;ۚ�cহ>I��D/���?I���?����?!&��7-���� W�j�k��O�:������?�(O(��-���O*�D��Le��{%��	oq���A��fn��	DÔ(����������ߟhɰiM؟��̹S��E����=g��q	e�	�M���?�����?��t�̠ڶ���1"d��Gb� c���;tl�vA�>����?I��?��C��$�Ӽiu��'�(Xe%O�7
D� *��ovX�jfӬ�D�OB��٢A"�I,�tԀ�f
�VW:p��!T-^��6��O����O4��o�2��O��d�O0�d����p��ޢ L��C"����ъ�LM\����I�n�$��o6�~����!�b�Rg�W�K�H+�"�֦q�	��q��Ɵ��I���I�?%��5����}�0�o4f�±+Ƽ!O���'��n\�Oǈ8c�y���ެQ!X���O�{�����M[sT�*a�v�'.r�'���O���'q�h��o,�k�
�-*��beـE
6m�8LR���j�	ӟ����)"C����M��0��48 ����M#����$�r�Hʓ���Oh��O߸X��*��ɮ���`�`
�yr�J�����O��	]mhQ���ܠkp�H١�Y2U*�6��Ohyr'M�<	U?U��\�	Z�ԡ�!��-� �3l+4�XK<��W~R�'pB�'��	�L/��0%��uML��"L_3%��坣�ē�?9����?1���FIk�$	�-�P�Ū��f�y�N�p��?����?�)O��J���|"6J�7�>��	B �v88�'�v}��'q��|��'pqOvd��nM�#���$�,l(p ]���	���Ixy2 �;k��୓�jP(M�ri��X�����NM����Ij��ڟ��	D^.b��wH@=s6��E�r�lk�-y�r���O�ʓr��{P?E�	���%�J8��I�x̅"� AW�ᩪO*��O8��e�<������32��(�T �tR0J��Mk.O~dH��F¦m�������?1S�O�.�#}�%��I�� X8 `�"?�v�'�""Z�yb�|���_<O��	B�A�+xn�(S	p:�����C~�6m�O:�$�O��ɐ[}bY����(R�-�e'= �u�P$M�M����<�I>��4�'�H��qϋ�f�q�D�a��E0��cӶ���O��$:;#�x�'f�	�H�m��b�aB�OsX�0���#XL��l�@�	�f4��)����?����N�s��X|�	��B�*î�cŲi/��دcf4����O�ʓ�?�1~L�)*&����0�5'W-{�R��'�8�{�'���'���'H�[�����	!0��0˖�§&Eh��vJ�`?���O(��?y+O*���O~��Gh`,�e�H�_餕��n��[�ʕ��7O���?����?!���?��'ܺ��T�A�J\�aP��)�"16�]-�M�.O���*�D�O��D�F���Q3�iR|8JG�&>����Qeيpzf1��OH���O����<9���.;�O���g[�Dt0)�sd���\���b�>���O��5�$�,~�M`�F7>�����2��7��O���O���2;]��'�?���r�,�%+B����so"����?�'��'$y��������[<W���"C�n=�#%N�M��Z�`3a���M��Q?U�	�?��O`PRw썭L�I���D�F���DŦ��	柄 ��*�S�k����/��S̺�۰��87	��n�y2�ߴ�?����?���k�O|��'�'8��scO6�pM��k��A��C(���OZ�1��Q��BE�I#mӒm�1�ٌp�DU���l�x���M�O|0��� �.$�eɂ~��~�%7�$Av�-���`1?�R��CSjc8��`�+4��S���B\U���<�b;+���FXF;����eA�G�zX:R�W�C��h�2�\J>�ڄ+��5U�u�2g�e�a�F b��ꃠ��W���y3e�,��3�D.��c6+������-��?	��?	��y�N�	��?��υ�?��u���NX�i˂Y@,9�0�'Y��(/O� �𹤈�%c_��ʂ�N3` "��'΄���?q�j�7A�8��6
����ߖ��䓗?���������0V~�Y#�O�B������	�5y!�"�
=��$K�4�<�4h��b�D|}�Z��ӷn�����O$�'9y�䁅'��]����J��2Df���?Y���?)���w�iy�!�9eefj����ID�pp��0FϠ���ڂ�Q�l��m��;2��D"��v�|-'>�����Lr�{��>0�$�Cc9ʓ87�Y������R��Fe1^4���,I��dj��<a�[20�JFdL/�fl�TaPYl ���I��T���`S�ER�$��e��*�ND�l\��15�i���'���B�L���џ ���^���׼�`��7��)��'�7O��BÏ:}*��c>�@�=�y�2�x��\2���� (�0��=0�,��>E��=krX���@]��E�:5j�æ�%�?��y���'�$�cSL\�� ����eu )s�'��KgDSH���V�C 5g����J���)X*��W��0O6a�G叔|%��$�O~a���MW����M����?ф�9~�w�`�Y��C~	�CD�5,Z�Y���O�}�W�(+�K�d؃������xHZ%��+r���AQ�
�4��5b�8S��8∠�ޟў ���B�.��	c�ҮTOv�+�䧟h�`D�O��8�����42���ӵi�T ��˓�3,!�/+N@ap��~��6�R�3 �Ezʟ��dE��iջi(���뎛w�F��� ��H)2�',2�'T���$�'��4�qA#��YL�1��ʗEv�i4� 
38�$�EϾ��=<O���gU�r�X��E�jtC�bY�.<���֜jL�l�I*<O���'F�虹x��XZ��?q�f�PDj��yR^�cT<�p�� hgU����yb-�6}̍2���h�I�!�y"(#�I�N����4�?)���򩜅"�-14# �(��а���u��yJ ��O�$�O
�P��Ҿ=�е0�'M�ԾL��|r���+@�ވ AFE�F�6ك��j�'�b5K��ѫw잨	R��q��Oft�oW�=�F|b��4y�� ��N">U��'��'��S>&�{E�����I�M�57B����z�S��yO� �f���dT�SKX17���0>�u�x�J�$3�h�5�Q<�N�8Q-��yR��2yQ7��Op���|:����?q���?��U#<x�ِ$
.�Q���Cւ�� AZ�:/2���>�O1���ș�<x���55���b`P!" (���G%��;qKI}���'1�i���Vc��H����)B�-K��J|����O�	*�S�#zЁ�ph�tV2�"�"O�� `��/� 4�(4A�Ah��	��HO�ӹL�>��Y�U�J$R���eO���I��JE��zh���� �	�,Z_wV�w+u��ܭDrҡ`AC��Z���'����P��W���t�!O�5����#7V( �f ��p���>f_a|Ң6�24x�e�	;��gC#�~����?a�����?)����$S�h���
�\��e��,V!�ě� 8�1�<s��p����B�Dzʟ�˓]�`@���i����`_�v�1���B��1yG�'FB�'_¬�v���'4�ډx�Z�ig�u��ȩP�Q�*���H�#�.Q{��'̜īG�G/��lH&e4h�$P3
�|Xĥ�p>��a�ǟl�I�Zc��Y�MD--p4�+�,R45�I̖۟'���?Q
Ĩ_*R��� �ɞ?}lZ8sg�1D���׬�N,&|��k@�}����mr���O�˓g���'�i��'y�4w��A�hP�q��1��H��3�Q؟0�	���#��)��9@��Y�F��	��S��%�[�21����?b�D�FBP�(O����#��l�2���$�'�O�TTP�F�A �"��ԏx��#��<b�r�'���'p�S&�h a V���*�fi�T��IL�S��yBʕ��5���"i�p\�l���0>ir�x�)��'.p8+&(T�.F��ۧO��yR��%{�@7�Od�ķ|�ꌗ�?!���?IB��E,uB��X#���̒�,��0�RD_/SΕ�΍��*��c>�
�GP�ͱ�h��K>�]��C�8sw��]�� �e��7ל��)���`����n=���Ċ@~l�u�E�7Ȯ����2���'�R�3�YXe�J�Գ~܈��'Q2�'<ޠ�dI�J`s�&�"�ح;����D�����#w'N@Z�N����01�F���B�	�`���x%��TJ*��/T!u�C��rɺ�"(�2K���)
�C�)� t��È
$,�l��c[�{�~��v"ODh���/�v�а��>�!"O0� K$��HBu�3М��"O�� �C	���3
�d�T�U"Oh�3��.|�pp,!�8[4CV�y"��`�~�J�� �zaP%C]��y��դsn�a��BC���ӭŔ�yr�C=}ɸ��V5
} A��*̊�yr#]d!t
�/��}�j�S����y�m\�� 1o�*l�j@ģY8�y��ĝ@b��E�N8Z�m�#k@�y��Bݺ8I���b��%�'CM��yRO�FG�k��ʍ"O~�y�$��y� �0x��Ds���9���˦Eݼ�y��Տ�Q[4*�>A���8�E�	�y/уaX���ș#96	1A��y�e��"$2��v�ۉ?�lXJ@OI�y��K���]��j�_'�l��D�yRe�2nT���eV(a�T%+�M�y�X�E�(I�!��g"�pp	��y�$�M� ��I�E"0Þ��y#����0�+ː=�d�k7��y�؍0�eS3�	I�8�+t�Q��y"*;Q��9{��	<H�~�9�H��y2��GM:��Blơ����R��yi�؉�VB����xk8�~�FԕR:��|��)�`ĉ�P%��{ 6���ӐMQ!�P�s8j(ʵ
��^�� �FU0{��	!5h$Cf��$~�x��Ҥ)��P�l�N��b�lR�0?A��X6l3�l��)T��l� >?ntÃ&�97G���"��s�Ew�<�s �W�}��G|bH�9&�)�g&�%��OL��`� ��I�R�(��( �'���� hz���u��&�"9
�':�-�"�ۈ�ܧO?���.I��3��:{�rXч�4D���`�[�{�՚ M�1�H�3 �6?��	�'����'?ySk6y��'�����bA�Vu�T���>Dt+�UU<�f��"#OJq�$�ف�d��g�1��pvT��j!�X�}㎰�H<�B'	Pm�n�:"EU�EԢ<!vL�V�' 2iip��q�'-�B��m6`ّ �S_V���F$�KybO$�|XC���{����.|����*�rp�%ȇ��䋨U=�Uۋ{J|�K�<���92�	��^�bp��h��,�ey��|b��f�~mx���'�$����Ǿs�r5�rJ[z����N<i@턖ntr�����Z��s�AN��~£M���=cr�Y/� ��^ަ	8FhA�'�n!A7�'w���ZcY�\pP�K�p<�\��o� ���M�%GE�u
�K�\�������g��oޑX���.��@�g��&~�ˇI>�@�lt��z�@�p�_<����VE4rd��-�?�2$ YHT���f�d��%�2�p
h�'�H��U�ޑ��a� DkF� �Ί�n�8�(VA�>Y7�7���I���d������TC.R�5xn�(��U���ǭr��mJ��I��ổ��;�DU� �|�(Ӓ�����ӒC���w%���݉���.yd�'�R�I4>p���a�7�����$�8�x����)��}����=��G�(;.hp�F$̵|�^�7(?�9��Oo.h����4j�μ�`DZ<������aZm�ۓ^VL��B�K/K�y�d��wN\�!*P;m��E����C�֖Y��'FL�#"@�M��솪^�6؊���Z:P�ǂVB8�<��+Ǎ[<H�D�+��,����D����c��J�(�-��� e1r��>A�)���I�)�i�'  �ǂ�b���QO?|���O�����$z�"�� @tX1�F�|��h��'\}e�Y*�!�pj,�Ģ�$O��y������њ��䞑.̹:��ƭ5lT�3�4��9�Ɍ�C�j�XG�V7~[�H��q�h��ϻ_�2L�p�ϻ�liQ�ޘ(�|)��LG����ɏI6|� ����֌Y��]0�	�Oh�顉}r�:$�he��KS?�d��<i�×�G���R�ר<�$�E!M�F�|�x@"j�z��W@X(4Ö�C$���֬Ɗx$�A)]���� eB�$�OB%)����<Q�(� ����0(�>ك  �$YFNX���.���*���%Iˌ��v��諂��66l}ҰĨ>i�HN70�h����D�@�n<A�J��6���R�����'���'T��
i���)`�ui��OԖ$�E���v�R�"U*�" 1z۴d08��S�K,ZdD2��;*˒�� nlgkޘw����U��>a�� ��ibl���?R4�}��$j�����Ǟ�����e��������c��p����Ή�7Ȭ rA�T�'{̅)s�e��[Ԑ��ӊ	:�m�4�N�e���Ȍ8����Q϶c��Ӻ��34��%i��AٮPgp�����4P؄8PFI$�b	�'�����.ԡr�"8�C(��p�b���e�6% G��9������j?�7) ;v�.�C�O�(�5Jɞ	�ذ�>�� �|��lx�m�*C!�<�p�ɋ�D̹M����ܐw�2�҇�`�yqWA�%
�6���EԸo�de;A-n�\�`�h�D��b�	�x��TRuV�`�پ9�m�p+�&��I�=�r��ش���C�7A����O6����P�r���v-�c�^-)����+�[d����c�?{ujHs��|�#GTu�R��1ր:�X�s`ϛ�}�T� �=Y�`�'��ޟȚ�5R��5^�8��Eg�f�J�2!@
~8�j��:e���ɷI�R����@#m��(A�7%�}���r���7�I	A��)E�y�<�I�?ѐ�-iR�ە��32$��X)M�
�������6-.� e�E9�RblW�b��k��)"���� eFvT�#�?ma� �EB���vO}�t��HU�A ,��Ǝ �-�j]���OT� �S8/daض�ƅ}��t���T>��g`U0X�|��%)�>�X�P��9�V�!�W���7�e���������y*�B-�i�	W�[�.j�Q�R\7f�hp�w Y�0�d��T>��2��.LX���ҟx)�O�:)i� ��ڰ	�l}�g��Ҧi�%L�y2���O~,<YV�5�����S��?��5����F�*b��9  �y)�?�D� �ѽC  ��	�'O�%�w鞗c�Шb�Ux��J��Ɋ,I�\���Ht*��BsO>l"��ɥ\`��Q�4s�$�K;;�*]��q�@��',�)���L��dh7��x(l=���Yp��� G]�6c,ъ���#
��(�=�O3���C(h�<y�M�	m>�-2�"OH� ��$BqX%=1��%���TI@:�C�{*��9�"Z:�JlI6e{��aCe�KTZ�a���k5t��t&4�Ot��p.8v�V�)@Lϱ@��kǋ[5^O���rbc�	���6<�T��,l�6�+DD?�c`j�D�F���U�/�F{r��ZqPq���+���B�ӫ�~��֍,����E����)U�*{h��@���0?��zs��ɴ+DTh����ޟh�3;BuB�.P}�`��!�|�DŨ;��B�O'È��c����y2�Zw�NL(�f�RO ESG��0ê�r���d�S�T"�,[$����H)~���PrY(lK�C{�ڴ@]�=n�}BM�}��"��
D�Pṡ� @i|$ b̙,<��[Z,��W"bF�� ī*t��h%��H֮�yg-ܮu�N��7ړ�ZHA�#��+��X	�c�S� �w݌�h�(޸j\U�k	�p��H�v⌅�ɐ ���a.�Y������\������^f"���IM�+�Mˡ�ϰ@�qO�S3ut�y�U
��u��XQAQ�S��ч�դ�#5jכr�P\�ŮE�T���1UE#v�ʧwe~����M�8)~���'�F����e�����*�Y(�j��X*Sd?M�H�Y��E�V�f����D�]~�L �'J^ui�bV�^<J���O�$pH�[���^#0M�PR���2c�Y�5�C-C�ў�� \3v�a8��H	�|�Tà��D˃��Y1�.@�kh��$� 4<9�Ti*�O<���&y��8�DM�3f�â�'O�m��K�c���8wi�l*=��{*��]a�M�{�$ ��H/x#�d$/D���1��(zʾ�3t Z�+9R�(��]C�����T>}c��V�r�:Uן�իM+~ (AEV�?�� 7���=ڵ�	�R�dd�	h�)�DfX%�y%R!QD"H(RA>*�j�!ES5�yB,��bu塦��0Z�4Tq-B�?�g�(to�=��I̹v�Py�С �N��&�x�ԩ�@��ȳ[ĝi��?u@Q�O�=�!��$��E�L�2~�x��!͓\r�\B6�'���+�|���9�4�h�Sn����!S�,Fp���'l3�ت-�2��f���4�}����G��P��1ɰ�(�B�xee/�I��^X��A�B����D@�'Z�hr�P�b���h���E�ɳF�J5G|r�A�&��ܚ�`�^y��'0R���m���4�%tH�@x�a���r��-��\@��4�QR`i�xbhSf]�q@�Æ�x�ݘk0����ħ51�@EY8��Vf�����u	>��`nF�s�n���`L(��#�Q̧`4x3 M0#j.�Z�j5��5�ŋVGZT�t�x]+��� ���bL݅�V,B#�':���!/��YPC	0Y`l�Յ�J2�ɢZʀ� gc��n�ay""�1H���H�o��'~�r�,��b<��j��7hĨS�B8QH#�?qQ���0:��W��4�BOҷOt4����L�V�*����'|$��U�M�R�:��ୃ��W�w���wa��s pP�ڟdzs�˫0�Vy�5�>�{��˧�Ώ�hx�B*P�F���	�i8���Sd'��k02�
d�V�?j���F��+w���'T(�/O���S(�r���"H�B��(CL�� �9#���ÓJ?F`Vg/�ɂ}*�L��O[�m�&R]���ɔO�����6) �ӑ�'�D}��)�X�P��2̓	��d��O��@1m�Q�`�'��>ɆŁ��� |i�d+�"]rp�;Yhp̇��Px'V�C8lء�Ύ� wJ��"�&�b��O��q_��e�56�,�I�X�3]�h&gQ;�t��g0sh C����%�R�_�
��5r��Z�L�#�<IR��N�h���Dӊ��P�B�B�tX*��d�b�h<0��ː5'�Q��ӏjtaxB�!e܆�;u�R� �nt�5�'E<a����F(����G�v��'����e��*`8py�dn8�\�Q͌"h�̕�u���� ��K5?)��B��v(B"g��o�:� ŏ�<,O��bnO�4�N- VIQ�/��չDJ:��E�ēcq���/��f����0T�:!8o�?t5rY)���|�P}�yh�'O�0�C�����6�����(���A˅e<�� �S�i�e퉁Sd���H8�$�'��Ӣ�-&R@��,щ@s�����mz��$���I�4H�Љ�o�5	1$p�
/O��C&�^<�H�'�ӭ0�TM������[�hhԒ���I�Vqqg��H�ԫ��VI��l�pe%<O�I�r�X�{�,T���h�Ś�h'�Ļ��R%�(��A��*�,H�t�@�J�UX�T�f�O̘��pF�<X��`�9�8`s�OĘR#_�1�f��ֈ�V�*�9WK�	u�r��o^9N���h/OT���\���bEpgj�]ڒ�R��Y"]���ΊF����6�V5�$�/-��u����J!�9�3��-7=�@�1	n���F��9�
�q�O4|�t����*�d8�7�0���,T��1O�3�v))FO}��H���N�(R �g
�'���PT�~*wF����tA�,C͙�lQx}M�Kj�d�`�Tx�8�6��qҝ�K�3��Z���/s|�#(͹>h�%X4���5���?U��4���n��5 ��2��S9���5��!�yB�м>��]#��P(2��
0
&� ``N��&!�(�n8E�\�3�&&^<S�띚A���2#S�g��ɬ�z�K����WOr)G뀄C�p<{3'�t���� #��q4I��I1s�0��WF����ya-�%Nu�"=�ǯ���p�i��.�ӿ3>E�aQ�k��l��┷}��B䉄kJ�J��U�7��`Y�Gιw�7MY�$��v�
;hC�)��튡�GR�$C� &!sA"#:D���p�Z�P�"cMw�6Yb��>���6]�ҙI2�YX�̣�ɖ�d�`��v٢����6�O�S�.|d��ۙ�jYXc�R{A�reSːx�k��&ܨ�#$ӄl�����`�F|bk��"̈�$2�Ӊ~���q �~ ��R�T=~>�C䉯<��D�T.;E�X�3�B��G5�C�ɖ.�<2�'� 8�X�#,SZ�B�ə[*�S�,�%GG�M;%Q��B�t͌��0	R5d���ҥ�T7D�NB�/]\��f-Y�#\���Q�M:y�VC��%y���	Qrj5���U�0@�C�ɰ\K�l0���U�t� S�ݥJ��C�ɚ�l\3Ӫ��d��0!""L�C䉌�e��L�T�Ҝ1��r�C�ɵT����)էQ7�PJs��4z�bC�/�����N�M^�!�Q @C�I;�DS����B���O"O3dC�Ƀ_$����o6��"��X�B�ɢ\�Y)��
 P$y�K�w��B�I�o����L�(��1��
�'�B�I�*�b�+B�WP�����j�t��B�I
d���:�'�$p`��+g�B�	�I8��`�Ҩ%������ߤY��C�I7M�H="����N���/a*�C��6m1�C���6x(�y7�R�(XC�	�Sf9I��]�}hy{fA�~K C�ɣ R����J.��2��6�B��S*�����Л��$�B��
�>�0��A�1��1!O�:FB��AQ�pHB�)F��PGż;B��<j�ỷA���	8��Ke
B�	 za*5�$��Y�1Rӂ�&!��C�i�jœ�j�2(���*�n���C�	�>�B����W+ir���H�\C䉰0,��!6fǌWh� N���� <�v`S>M��L�ɗ�_��S"O�m��(9�l�8�-�;�Ҹ�"OH�q+.#ypN�U�8��T"O��h����	�n�Kg-�S�v��"O�13����Յn��A�G�V�W%!�D�1H�`��Չ
��<L�
%�!��y�R�CD-�%b���dl�87�!�d4Q6`xс�j�thUl�� �!�Jrs������C��KY$)�!�䚛/�TB�a�9x9r�Ĉ�/9!�$/w��`t-�),�X���#ק8%!�d��"�ҍɖkc��H�(Z!�D�}�,��IRh��˷ǟ�#!�F�G��X2��v?F�Is�8P*!�$�4��ԫ�H�%"8�<9@�ݑN!�d�eH�Q���(�^uJ��ʷ�!�$�:)�T�������A!j���!򄑟�|\��(	�.���ʷ��sW!�$И0��A"!�.o�
�:P��}:!�$3jZ�URC��&���7H���!�&�&$B�.ܲMl���#h��!�Ψ&l��t�1
e|@��[�C~!���.��喾L�h�RRo�5!�$�*��<��+�/gߐ��� O'^!���A{ae%�| x��*%!�d�.|��Z�)�����(&!�I4d����6d��8%E�5�!��]��*]��/!�����EY!��Gez[��&�\0;ЬR=OP!�dR+cU\-�΋9M����,�7}�!�S<J�r,�u-�@����H�!�$�0Ea��{��I��l8ƠؕK!��n��b=6H���t4!��ߑ~}�%���u̾�3͚'L�!�dD  ��\BG'T$:��!P�!�Q�!�$� J_�y���VBن��3��<!�DB�pA�p�Ń�pi1G�EO��E�'E;]��(Q�ʱ��-����y��Y�5e�t$gШ5��%���A��y��E�'����R�ĺ ���gŕ"�y���.�
�Ȅ{Sz�����y"���4�"���t� E��I/�yҬ�a.4c�$��5ű`i؍�yRH`3h*�^�/~�ш�/�yBZڲ���ݤ#����&@W�y��	�D��XPF�X���'J�J���%�� w��Б���;��2JM8"C��X{�+U E=5����&Ɗ�y��C�	m������	I��ܸ��I�-�nC�F���h��)=|�{7��n�.B�,Z_�2u��:Q�T�J3p5�C䉇�f�hu��/����E�$�
C�I:%�m�P��P�j�a�
1J�B�o�@�[�J�	i_����CA9F�C�
h�"$3�C=
r��0��	�&&�?i��X�0B�Ѓ|��@��ɐ:n&Q�ȓZdAb�>?��7#�T�q���u���3�.��T��U�I�ȓ~�=;GO}�ؤ����)|A��K�p`*t��b��Q)�"
L!�<�ד �� )5b/h�;��Ҍ!�`��"OXEH�4���
"P�L�LT*�"O�쫐L&��"6ꑐSOHu"O�8U��^����шեDD2�����Z�� n=��i��d���X(�>�;�"O6�)C��l�h�"[���y7"O�5�@%��Bh[�?��Ɋ�"On<�D�q�ѳ4�ߓa��e� "O��I�"��dd��������B"Ol���������bO۸	���"O�S��R�:��)�# �S�0�V"O��xeDN�q+�EӶ���W�jysT"O`�2�,{�ZPc��	<�$��"O��H��ح!s�;��+CV�P"O�IJ���4��ų�C�p(�Ia&"O�3焟9T� 4 ���-o�xj�"O&�©R�]����R 3"h�W"O<�r��[���&���4�z'"O��dԔ���1U
Ƅf���pE"O�i&	ؕ ~� ���%�L��"O,��uǐ�z���b1��.�>��7"O�L�w��#ưd	��I>k�(��t"OB@�� .�2Da�o��?"\i��"O��iϐ�&D��O�
L{�9d�'��'�Ifù �j�Z�N�8���'A||aǡ�*4z�K��R�>誈��'�F=��w���1�N�9Ll��'y�)�!��P.6@��ɘ45�8���'���Q�kTDA����Z�	�'DYk�/��ܨ��&�\9��'�8AXA�2���`!�Y�(�� H�'��\1�-<2�ֽ�P�Z�'�Fȑ�'˰��)Qr��iW���&�"!�'	&��@��9(R�k�cЙ�|���'�Θ��G8e��YY�À�c,lz�'jDZ�mJ�W*�Z��²	#8m��'Gv\J��N$�H#��/zOBr�'����n�R�W~���J�'�"(�7���E@���r$���
�'`�m��b�H��E��!�b��PI>q���	�1y@LpR��(��-�
6C�!�DԜ��)Z�%��r()�AN>!��{̝yɇ�
��"���~�!�ĉ� �����Z9|)
!��"�/$!���%yL�H�I��h�F��!�F
\؍���E,�U�HQ/��ȓK�ڝr��ԬSVl�D��1����U��D:�N�t^�sN��j(���r���W)ǜ{W�Q�
Ì� �ȓ GBe���."��@�W3 �A��~�
��"*kk�0jɕ	&���	��l�� L}��aD&� .�q��~�8j�Dشt!�1C�Y;,b�8�ȓ9�x�ۄ�7��y1.�}&Fم� R}��O��xA�m�(ưS�}�ȓl&�a{�B�}c�U)7h��y�FՄȓW��
5�	;@�L���i�+:�\I�ȓ=jx��g��7%�Y��]��Ψ�ȓ'O�P�6�5x��:2�	J�&x��Tb~u�%!%�4��m��##���ȓ�A�i�����IG Zʤ̈́�_�|�S��B�N"dЉ�G�9@�@0�ȓW�4p��
�=�Q-�n"����tIQ�ӟWXu�������a�Q�`OϽ'A�a!ւ: ���7�Es `� af� ��|�t��	԰\U�5#PnT�"��8<�ȓeSjر��`�~XK�(K<>܇�S�? j���ˊ�&��L�+T� �"O�LX����H=��+�o�8}� "O��Cw��?�����Z�SfJ��"O&}��Ĉ{���U�V�V�L�"O�t���B/1��9���2m'�%��"O��� �@3dVٴj�[{� �W"O}�2bY�+S��锩�g[�0:�"O��1ą-�l��F�%nh�kW"O�,EH�_���V�1/D�kw"O�i��m�460 �!wt��r"O����˛��  )شVn��"O�|32b�jZX��Ȗ`�d}��"Oٓ5��2x6Zt���ςY���q�"OTp�!�ժZ0+��)-�Dģ"O��%���	��/��P�"O�l�R<x���+�̀D�P�j"O��[ъ��l����C�	���"O�-
BNӉ!Xd���͓*��p�"O��s���*J����`h�4Ʋ�:�"O�Ȫ��V9�0�1VF})%"O ��`����9[L��]pI0"O�T�2
���3%�	��d�"OLd�C�_�-I7*S(W��iQ"O�a��D�.��-p0�H�U1�"OH[pB�/.t��H�M�\}CE"OL���e�}e�R��[
k-$�A"O�x ���%^�����^
�x5"O4%�E
4y�:�pF��
S\Hc�"O��h�.
�e4-
D���Y�0M�"O�IV��iDNE�u#����"O��!�˿g�����5d�V\J�"O�, �+^�S"`�!��݌X���|B�)�Ӭ,�#�I׭U�F�#Ō��C��4'"�(QQ�$X�|0�Ae�C�I�"^���rŀ�t�v�@�-GK�HC䉵\��D�pᚭf�L@&F��lB�ɰ-��9���?O�8�I�,Ĉ�XB�	hJ�la���,��|#3����"B�Ci��[6	P%_B��""C�jrZC�Ɏ+
�5��bԚ:�,j���	iP,C�	6��T#�*J�x��h� ��!��C�I2F/���v@�1F��T�ɒ.��B�ɩ���T��:O��p��(x0\C�I�$��sR�J7rRt�b�+±�0C�	c��m�р�� Mq!f�V��C�Is*��x5�C�x8���ǚ>j��C�I�fP��k�i�L��(�C��5.���+` �4��W�(��C�C�8L���JC���ť��J�C�I���-��,X�?}�8��L�q��C��2ƕ���6v����P�g�vC�	�,�^��4���
���{�$]nC�I6sj(,� ��	enL��'��@��C��;��P�n:m�$ Ô��P�bC�	>	�� �iN�k��dÖ/N�0��B�$'޽�AR7"��y��A�`��B�	�?����(Qp���ǟ�g�B�+E,�y`����[\`�I���C�I)������)}�"\Q��2Q �B�	G2`��OV
(P�0c0��.=C�I8 ��X��k�cDePc�;7�6C�IsSf]#&g��&�.���矩g�PB��
r]^�[��Z|�,uh��I�C�� H��� O xI�p��i�,Y�|C�)� �ڢ��7zk�a��r[�3"O�I�§B=~�JP��ˠ?�%�"O�=B�L�
_���Z��O4��8H�"O���1,Р\��C�B]�zz���D"O�%xS�S�m�6k%B�0_dԁ�"Oj�Vl� �X� �+�o?���D"O�	��;	B�x�ǯa% �@�"O�t�F }�\t��c*"�}u"O�E�c�,tn��7b(&H�"O���A�T�����dB�k�XA��"O��qҊj ��W��z�2�"O����m��*B���H�R�*���"OTh ��0q��M � �a�8���"O� �5�]l~`-`@�%n�6��4"O���D�<?�d��$��Xp��0�"O&�c�OŁ�\ău��ad\�2�"O"A�卅?�)y!LT�>����"OX��̑3F$�36%�Q��i"O� �f@�;vzBI���-
�(�"O�Av�I#fPP���A��Ha�"O��BT�"/�`l
a�;�d�:#"O2Ԁc�V"%�N<)4�p~2m��"O&-����.p���&gܖhv*���"OfaQ��O%(���YAij��0"OE� �˿dtlh6���0��"O*q�TB{��x�F�&�����"O��2�G�D߀q0���In䂵"O\Y���>��M��,Qd��+w"OV0���ۭR���`?f0�d�q"O1QM�~��j#�%D%Ft��"O���ԡ�.ʊ���GT�J��8�"OL��Pj�!I�*t�1yN^8��"O(EJ��^1hj̍"Ck�.l��M��"O����c�J����mv�2"O�Z.S2+/��2�F7F �"OR�z���47��(�E=$��D"O��c�� ���q!�#uVQ�"O��BP�Ѡ%l���^#_k�%ZU"O��b$E�e� � -2 CRP[�"O8����"E��=���W h0T��"ORlpפ���dS!+��s̵�"OͣD�R�y��ѻT£�H�"O���'�E�Q�P]�cJ��}�*0KP"O���g�-� R�H����3`6D��B�˳*�F(V�O�}���cTj7D�,���@���ӱ���ᑔK5D�h��R�|��4��g��	�H���3D��t��+(ՠ�*�#���A�G�2D��t	E"&۰h'Oۦ3���`E�$D��
��2ޜLp�פt^MPp�$D���0Ȇ:����WH�F��𘕢!D�Xa���h�����N�4.yY�v--D��1� &��ti�D2a��5D� i��ԏۀ�����Fؚ�'D���n޻�r�
��J�:���G3D�TIM�T+�q�e��1t���'&D�$I M�)|��!ʇ�p&`U��,/D���O؞Q� ��ר� e:�o(D��a���DZ�Ke��6>���v�"D�,���HL�ը��L�49~��VC D� ��"B-T1��r��4d�:l`->D�����.T�1��$H����s%<D�0{W�Z�p3�;��*��4�Qh,D�,�c������J4ayP�(D�� v���I�{���~����"O-�5,��Pa�yq����h�ؔ+�"O�	m��7lX+ n��'��
2N&D��Y3��8�ʡI֊�<a��z��8D��ã@��Mfh���kU����1D���p�r�3Q�Q|h���1D�pa�iǅ
D��(�%̻,f,5B�./D�� Q�	@�s#�^�\�R�7D�l�+P!)��љ�,Q$f'�qBQ�4D�cЎz���b�Aez}�W`0D��[���32`R�*�W�>W�1�y�dɵEI\�qF��<g��yPt#X��yr���J=�h��j�(�����lA��yR�)1)�(�U�K�v��8դ�?�yb�G[��bȖ�uްQC'M�y���>\۠��b�0o*�
��?�Py҈]�?vRYAڌt��(ӇӬ�y2���t�!w�@�T+X���G��y�i�%��8r�I1UgRt�q�P�y���m�й@�P0O��E�ܕ�y�h�).�8���i��|�fԹp��8�y��ƥ�$��+Ht�&8����<�y�h��P%p$�DE Z��Y1(Q%�y�+�8��X`#�J���x����y���5)��āǪG��ՊW���y�F�r�\	�1��@��!Ǉ_-�y_�D'��vW"7y�%����yÔqME���.��a�Vf��yBH�h0X���X5���M��y�M2�x�8ǎG+^0�|A�Ć��y��]m@U�E�K�R�V�C�D	�yB"�z� ����ؚ�W!�y"�H�^�9kt��U�T ��Z6�yNޓy��K�+�M�d��rɕ�yb�.y�.����)H[*i�ҩ���yR��*q�V�톇*�p�9�,��y�/���-�wUr�d�4�X2�y�"�5g�QH�9r!l��2ϙ��y��
�d��)c��~+$q�w���y�������3,�:M��������y"�A�8-�a���zm�`r�e��y2���-Y8�"�"�D|H$c����y�'�x��E�%[�՛�
�y���S�h�Z�dÇ�t��͂�yrnE�n\ڕ�A3
`���ٮ�y�8bV9zvbN�94
�pqi߱�yB��![�l;e��13xx	�o^?�y2��/Mo�#0Z����yr쌑w�����Ł\�Ԝ���K�yR+ĝ`B�I�O�:�!���4�ybA#�<y@1`^�vђ�aĜ=�y"aE�t�0x@G�Im�
Ÿ�l$�y��ǜ[�񬘛g2(�"�K�.�y� 9J�m�A"F�H06�D�؂�yR ŉTo��!5�@��q�$C���y�dƬ�\����9F�+a�$�yRgr����BѫL,�1jЇ�y��L0D�ʕ:��L�J�B�A�܉�yb���i}��jd@
�;�$E
1@_��y��7QOzai�?1\�������y���vPx�qk��y�*xS���y��9x����P�~�F�℈�4�y�N�Tp�I{v�x�U�t�A��y���������Ůo��){�-X1�y
� f��g�\�%�
�Q4�K�\��$"O(�e�f�Ȫ�� �z�Ơ��"O�I�Wi� ft,�c%@�]�,��"O:u��d�p��0%��|X�1"O<Ƞ�A=l��u7����G"O���h8I��h32�-�����"Om �,�8�j �&&QY�a""O�買�0+�yx��AG�t|[�"O*��A� 	�9���A�?<�"OH-ذAtS4(�h=�A�IM�<�!��>S^�x�S'��M��y���E�<�"Y�d&%;Я�!\Ͼ`�sG~�<��В& x!��[YR<�5t�<�ŋ\w���ę�<�����_��`�?i���OX�$+#`M^Y�X�A�"��q�!��L�#��	����x���*�!򄄁Yb�Ŋt�׺~����&`���!�dW v�p�(��d�ݟ&"!�Ě�l��W�K�bĀ�����-!��\r��ɷxb����Z�O+t"���dOw��4h "O>�CD��JR�I`����Z�s�"O,0XVj�54�����V!�|���"O�h��O�.��с����� �"OP�!dB���iGb�6 ��!�"OL�ajU<���k	x�JI�"O�����X1^�(R�\�W���Q�In�O'����@d2�8����j�����'&,�Ph�z��3���5�ڴ�J>1�|�����)-n	���G�$�P ��4�R����1cg�,��*�a��kCp�7���V�DA`��7����#"x,�G	�6ɸyd�7q��d�ȓEoPD5�]'B��mY���L�&�܄��<4�V��2,��(��H:#Ȅ�`QP���$�	�l'���[:TJȠ�Ԉ@P�C䉷�~�����=fёB���8�2C�ɸ �����#n���G��P<C��9O��恌m�� �T�_<�,C䉏�.�(% [>Դ�st��1z�@C�ɓ[�Z5�+E��xa�0Z}&�lD{���
BoX�$���6��+.�y�Dt	�C��Eh��A���Py��*z��y��ɋu�Ԍp��F�<u�ݷw�����JD�D��$jB�<�팮q���x��u4�`���F�<��D�6K���d�3\����N�g�<A�ܨ
 ���G05oJ92�A{�Ii���O
h�AP��iX0�!5�L7)�N)
�'V`�aJI;@A�q"ďk����'w�p���>*�H��J���hY�''���E̶	�����)�7|�x��' dz���g<�E��{�8L{
�'0��&ղ��%�눦v�ni2
�'��+bD�
e��b/�$|{X�B	�'����肺+��JЩF��TP8�"O���i�+_z�=��+f�:ahp"O�D"W�ɸe՘���l���1"O]��Ȟ�F�jL�R��7⚰R�"O����d�D������v͠4�4"O��az�"p���� �uQ�"O
�xR�9p������$!?�IP Q��G{��i��<4G�r�0�u��r)��V���RgM�>Cx�Y3 U��M)f�6D�� < `iƵg� �J�f�(�0�"OR��F$կC :TK����	��"O�гc�JE�}�M@�]3���"O:�K��B���I��K
p��Y�"Ox�Yq끽[4��J�iہ%b.��c�$#<O0YRӪM+~!���R,h���X0�=D��q $A4kwl��1U��}c`B�O���hOq�d1��A���4��9 ��u��"O�]�"-ڨ��ir$œO�2i�2"O�r�ślh��Q�A(��`A�"O`�r�JͰ-���rw��$�ܠ"�"Of=x�@�2tW�p3B%W�����/LO\D��D%/w����v�A"O���f�����@�
jvA"O������ߤ��ՍD[�а�"O�h�QC� �Ȩ�B\NQ�x��"O�@�oL����T�X�/N��(q"OL���"ޤݢ��@�3&t�:�"O"PRVD`����/��
�T8U"O�h�&��Xk@��%n֝V�:)jf"O,5��Jʥ#�
NA�IЖ4��"O�m�7BM�>�r+�S���p�"O��PW!9��y۷��l�Й��"O �k�
�d �q�߬2�!"O�E�"��OE�!21�d�$�"O����)=(�fpI6*��^��`ٶ"OR*1�Jv�t²��=Yp�q3�"O�

 �-є=S��A���4��"O0��b��%D��S�R����"O\�xGEN7i
�3����*X�e;T"O>H�'@����*:U~�R�"O���p�C����K�˕L�k�"O�ˣ�Q�f:��@�mL6u�b���"O�Pxt�L"=`�8�K��
2б�d"O`����+�@��jJ��a�"OT��a�7c����cS�o��Pd"O��q�
S��0 �ْ4��+�"Oܙc7 �2P�Q�w�5�2"O(,�'�`��)�c�I r'N�RD"O�`{�D�K� y�5ϓ�v��p""O�5�@<B Ȱ�4�U�N��Hw"Of��"�
 o����l�7�v�7"ON�c��(�ڸ�DE����w"O��� "	�:@ZI �E�(�� ��"O�Xd� dL[V`�,i���"OL����9 �r�B����mF�p�"O�ȳ�KD& �(X����Z�4��C"O�9 l@=a��B�FޘFf����"O<��4n�	a,D+D�G`���"O������-WPY�ޣW���g"Ox �O�"
U�&�D����"O<U�QM�Fa���/��æ"O�Г&눃S.(���o��7�TU�e"OF�q�EC�7��p0�ˏB��@�"O��K�D���������k~�Y��"O��H2M���Q�)�����"O����D�����b�I-h]J��"O��ò��3B�x�ʁ�*�\��r"O4L�4i�(��x�UG�m��5�"OT,j��N�HYthI!�A�Ux\��"O�IxU�B�b���&��a���"O^�k�i��g�\!�!��R����"O�EJT��\쩓�N�E56tj�"O� 6̌�7�6i�qm�!-`tق"O� <�9@"C�G�����]9��"O��d��"�̹��ް"uBu0Q"O�tyS��]?fx�#�3L�"O�E���_tDrX"�6f��!��"O� SB��$���;B o��Ż�"O�kO�pt��.J/�m���"O�)�"�Ma���cn@�eb��q"O�iQg������%(_w��`"OI`���$-�68���Fr��"OH9胋�:;��+�]<Sp�e2`"O�Á��Y�Z̑�©e�T�"O�ɘ��haU��-_(�i��*_\!�d��4,���de�{E`%���F�C]!�d�CQ��ke���G��q!S-ǠNY!�dD!=NJ�Q�$_Ӟ� .���Py�(��s�db%��	w����֫f�<a6e�f��ث��9D&�ġ�χh�<a�̜$S�p0�޷C�|8c1�J�<6Qe ���*ʋ !��
s�ZO�<1��V :��x�,�
Q�^ ���r�<QSjI{)�u�6���q���@cf�j�<�Cxή��)�H���[CM�i�<ёG���Lم��$�T��d�c�<�[���8#�
�l�LxP`�<	�Ӂ5��b����>Ԋ��!�^�<1R�F�Z�A�b�ʏd�0��rj�E�<a���\����EZ��L�Z�nRH�<��4Z�~5J��ߚ+����GA�<ɔ ��^U�<C���m��C���~�<�2B*��d���D:{HDm��J�e�<�����~9�u*�V�]!���c�<�Q혘Lq�=���+{�����c�_�<�aH8��Mq�)S%}\��`���[�<	W�J�b6�ct�ˠ!㈍�lM�<��eW?0��<�tL%%��H���`�<	��x�4L@��"?(�uD�_�<ѷ�Ϭ����JXF��Xcr�U�<�S!A)1*"�a���*-�4�ȓ+A��h@m�pS�4���/�f\��_<��볤��z��ĻF�үz�=�ȓirD���R� �1�M�&��̇�d��iխ�/'�pٱ6C��\V�e�ȓJ\ hj��cB�]A&bP�\�ȓ�����3X���@�j���ȓ����$'�4M@�Dh�kM�fJ5��w�R � �V�K��W%J��|�ȓ5BH!�e�&����[褆�DR� �&M�Rޭؔ�E�j<��n���Q�պ((勔M�6,��m�ȓc�k� �%����9.�F��ȓ>��X��%YiD��EQ�'���ȓ�4�)��Q����W��[�z��ȓbt�t �_|�H9�n]S`jX��*4��&�4*�MX�Ȅ8E�ŅƓ]�
�+���f����S �,�"O��آ�N�,�`��@T�gl��c"OL��O��D��dJÎ��%�	q"O,yp׏�XQ� BR�"7�����"O�|�HF�)v>- �J�=�� "O��w��%c<��uԴE�X=)"O|�*�����
(v*Hy����"O�!R�W�ƥ��o�,0}Ή�%"O8�bVdFe�u���5z4X��"O�U� ��-��H��V$=�2h�$"O� \!�OF4��}	 �d4�s"O$�dStZm��*�j *�t"O�z�e�nR�*&,����"Oj<�&�S�T.ZH���µP�&�)�"O�n�dy�╃h�2�h��P&F!�$�`H�Y1RnO1�d��"
O!򤐤2��y�%.��]RrBI��!��Vusѫ'E�1i|�h�A�|!�@:8Ԁ��
�?13�pٷ� 0\�!�d�T=��ّ��#A�RA�OU!��]�6a���aq�A�%ݰR�!��ǣ]`�Ag�oD�"�@��!��N�T�8�B��KZ|@�EN�.�!�Dڅ+��@���f>�����!�D�	S�(��Y�B��0M�N�!�D�!t�Z\�N��܌�1a�ͬ.z!�D �w.j��nȈQ�d�1}�!�dM�	����¡�,���!�L�n�!�$_$P~�$�fJT�� �'ҹe,!�Ɲ�p  �Pe�����3jm!�O�)B^�R�eԯG���f�I=N�!�$�
[/�)��H 7D ����I�!��d�v�1��83�G$�\�!�d�&�p1k0!_)}Tl�<G!�/\.� S6#�a�t�lT�,=!�N�<����GG�s�ꕴt)!�$�+b��h@�-C8�D�fHV7c2!�d˂Rxu�1�S.q�Nx"�LҽW(!���.�!x�	/#�)�%�ǀ#!���S%��"t͏/$h�g��e%!�I1}�<ܘ�G�f�i)���+(!�B�g*�Z/G�
��M��%�w!�άZ4��jW�o㎴���ߢ!�� �,C��2��Gָd˵��1.�!�D��o�&e����"d���	��T�!�����u��� Ri�l�!�dǦ&q8X86�|u�S鋉hZ!��+M�R]�&���a^���,mF!�d��
�X�ã[�{2��Q ߿5'!�ă�H�H]IT�P8?y�騱H��!�D�:wߔAf�B&4m$LsԦ�L�!�Q��ⱂ�OX�$0`�N�!��*B��:�aƎ[���Q�V?�!�dH%G����6��q޴��`���r�!�� 3q��$��>)�*��21T�!�D�QP^�4&�&&���t@�!��+' P���ܒ5��q�GJ5�!�D�:Y�2�,\��Jl0�i]1#�!�$_�� �#&�s6"ȑ�]�!�Z8eb�X��S?S#���F�N!�DR�)M�y2�IƝl>�9�t�Q>=!��,�M�#��@BL�)�tk�'����Y�dhB�ѫ��ɒ�'I6�����0�mE��*d��'M���LA��aAﲍ9�' `���`*�8���V�?�`q�
�'C@����n�K���2��p
�',lu�ݠ%u@�9`�&��+
�'k $Z�C� "�= G�@���8�	�'�@E
6Fi���3�i���
|B�'*��-	/Ql�0:�뛦B�H�'�|��"�vt��CJ}�h!
�'�DMY�CW�
D�1��qp0�	�'(F�k�o\|yҀ��e�Z���S�? ��BTI�4SNf);���s> �q"O��饴�6���y�@���ʽC�"O�����\?�J��GF
�l6�!F"O6�Qv�Z�`���XteŇ!jőG"ODh���/�m��]�]p��2"O��� ą	Q=}#蒋� 8�"O&<�Ș<*h-�%�
�}�
�9�"OZ+��\�0��MS`�׌%��Y�#"O�D����F
�8ƫ�B&���"O|"��O�w�9p��y�NA#�"OD�
0O�9m�̳gD��Fd.`�"O��@��-���r��xaJ��"Od%���9�R"ӂZ_<��R"Ot��uB�.�I�C/~�᳅"O4u��`E'����a�ij�Q "O�X�-X����3�%]���t"O�s@!�' ;��9f�ފZ|���"O�U�6k+c�rM�R��s=���"O��(p'T�`���Zf�k�d"O�*���d�����k��^%ΩQ"O4��V鐹X�(��F�'~����d"O֘"�H¤4m�"+MA���&"O�l���E� AB�&�V� A�"O�D'�I/���RG�]1���e"O��JF &2d`�炏ӊ���q�<�i��@��U���<�4ĂAL�Q�<yq�\%L���ض�*X��x7��J�<ARI�*��D����$��@���C�<	��Άu ��ۄ-W�$#b����	@�<q[�U�G�d�k��%�4��9���R���V��`���.�ȓ-+V@R!"�6*��8Qs!YW�rM��`r��q$5������6 ���۪5r��v�ӗ�"z}��L#��
F��F�� NW
yv��ȓ`"�9�N�_Z�`�P%>s4 ��u�|WbF 	+���� ۤ��ȓ��X��nS?̔ ��Ir]Ȥ��x���ǎ$���Y䯅km�ȓ0� �Á
�i��Ap���Y)�ȓxP:��ܸ0�bH�u�4I�ԇ�9Ly��@B<�S""�Tb�$��*���F�_�Dذ�c�K4�6��@y�
$�ҳt>�#E�3�4�ȓq�$h &D�m�䌩���~X��ȓ2*0���)�%3��K$��tO�̈́�\�<�"]�x�"Gڐ����N@H�<A�ZR�������U�h�p��@�<! �5N$4�&��6����GL�<A'��1B����AN�GƼm��f�<�`-��򁱗��4��A�o�a�<�d�	-N�yR��>V*�ɧZ�<9�Ą
{�X�ᙂ	�vQ!�@q�<9�H��F� U�sC �=`9Ï�T�<�W*\"_����`�C1�daQ�e�<��� Il	�S�5�tIy��a�<If���5�L�5f^LP��fD�<)�Ü���1T)�d��"��V�<Sn�N"�L�u�ӊg�,�ƨ�Z�<� ��J�Y��Ð�(T�<�d�� ~��1�jĈZ!�m�+I�<ٲLځ<Y��D 9nt0;��L�<A�hB�e��@9G�5[iܙz&�	I�<9nB��V�@��W�1��#DC�<� 2�� ܕQ��L��|�T�`t"OR`!'-W>8���r�O�b͓�"O�����>I h,��.,��4B�"O���a��6A�U���լ{t��"O�y�A��`��0UmW+<^ hI"OTe��M��[p��V6n�L�&"O�a�J�=h`�x��A�0]h�"OZ|S�Y�t^����]�2/���"O*�xX)n"�TlܔX�8(���{�<9�p��%��[*��#�^�<��Dݙ����Uf�i`�Tc�.Oq�<����P���W��	H�ꄆ�f�<ٵfK�S�P9ӀhIGr]�w��\�<�"F�~��L;P�XE$ �#�!�L�<9P	@�|������M9HU�Ad�b�<!!�ua�e�k��٩���`�R��S�P7�Jݔ���ĠbItY��\�ⴊ�!U%�Bܨ���b���@ᤤ���3� ,�d��R���ȓ^	V������8D��I\&:���ȓLv <Z��ڮ,���t�"wn������ ��B9~�8�&*lͪńȓ_'�ɓC/!8�Uȱ��=v.0��ȓ�0|��ɼ+M �#�J?-�����}L!q�@�GF̩����8�ި�ȓ8�5s� =~���%F�p�F̆ȓ�N8c�����Pv�Q��-���@�jE�X�krq����$(Ň��n�1�,"�h��fAB�Jt�ȓ)5�T��I
����m�[�bl�ȓ K�iЖ���U2���4�[�&ŅȓZO�4p)�����1���?F]tP�ȓjZ��t�1|��°�e��9��o"���C�v�4 �-`k�ńȓ'}P��aBF'W>��C��n�,�ȓQ�	�ɉ
{�9yB��g�ɇ�)��,K��V;h� P!��"��|��IRJ��ʎ��� 	o6Z����Hq�)²?.0z��1�)��k�ĠG
_C�h1* �؟
���ȓXx|* ��$W�t��!P�-
u�ȓ`�U�t��%�px�&.4���ȓ%
�بJL;0|~h0�e�*2n��]���J��ÿ���O$�|��ȓW�U����N��{�Nثn,����]g�u`�FC�P���{$O�rWvP�ȓaO����.�}H�����*w��y��^�E�tI>L�iu) 'e^ �ȓ��d�B,&�  	�._24h��T��!VDC#.�k$�'.�&q�ȓ:iJ��kKA��a���j!��ȓ,D ]�	��A9[3+�h��T�ȓ�Vx(��N�TS��2 �X�?��݇ȓS@�ZQk=#��P�	Se���ȓ:�~!�`/ǁ_c����4��7,�ݫRk��as�"�n�s6l��q�8�%Ă�:��=�R��Z�9��{wT��'�:3�@B'C���	�ȓzp���bV$=},�"���P
\�ȓ�^\)�
 f�lJ�(��E�����7Hݩ�� ޙRq�U=h FP��*�m��Qy4|R��ZNT�"O"��7 �d1c��+h��br"O6!�Cj�@�e��T����b"O� �]�`ɚ8E�A���\�����"O:�:�
�B&��s#�P��+�"O�t��&��I���:Ζ�q�"O�=aU�K�a�NR�����*�"O���!��`��FKN�\� q�"O�HR'	�Xn���A�	� Zf"O:I����N��M2EH΋K
UR"OڑI����f䉒��	�P ��"O�����;(�І �
&��"U"O�JQH�rڼP'B��1�|4!`"O0��� L8P��
�p�`$�1"O��x׌�U4" �؞r�:�r�"OX���//��08�l�*$���p�"O^��qa�8mÄ�t�V9��x�"O0�q2�/U^�����\(0��iK "O
��M��P���OQ!�}��"O�y�J�?��г�Ƃ��"O�=�v�Z<L�
F��/W 8qy�"O�!�2�ڽ����)�� M�؋�"Ov ��ˆu��qkaIC38VX���"O�T�G��^���ÓHȼK^n�"ONe[���6`�d�VHTfH�l��"OTcF��.WtI���&WH��"Ox1#$�*j�V%�!� �l8��)�"OX0Q$-�6rP�}�����"OV�hW�˃C�h�'b�<�5�d"O~墄2+���t!�5�L�"Oؐj�ɔ<�6ՠ�<	 �e�D"Of�Y�Dޜd�BP�ӢF�\��1"O0���MxV�|�K�y��R�"O�eY�D<?�Z���g��	LT�"O�E�� ޙ 踱�� ~)�Ē"Oe9�֛+���hΨ0�ԑ�"Om�K�?�R�Y���E.N27"O~�+Ac�,6��f�6ʺՂ"O^�	���7 ���6s�%�W"Od@+�]�g��t��*	>!Ȉ�6"O��DES�-'&���*��]��p`�"O0L�Ё�4��A�TCD�F���"O^e�-ʱ^�}�2c�+{�8B"O�prƃ��&M:p�G��oz`�`"O~�[S��
X��RL��P�"O�䑧q�<$���?a���z6"O<�C[�M��䃶���X-�"O��Ȥ,�U0N�s����%'T��'"O��tHڄ����/
7^	�Q��"OD����ņp)X$:��� bZy�7"O9k�U-B�`cF�������"O��	���NjU�&K5�N�C7"O��X�*�>w4x%���-�
�"OI �J�I�x�h�g�(�Խ��"O�1�g�7^��  �B|�l0"O2Ys�čNO
1�g&�U����"O��+фHV3�DkD���Z
�A"O�<�`gՐR���D؉�\H�"O�څ�,7�Q�-��y�RQ�'"Oִk�,W)���!�m�h��+�"On	� �i���X1�B(x���X�"O�Öh��)�&�|��`�"O�M�Ǉ�榙rD�;k�n��"O��0$̧c $q�)� ���r�"O����$V��1��Ċ�^]�S"Oڈ�ul�k�X�B\
I�L[�"O�Q���W�02j�PW�_� �B"O� �Ŏןr�L1�J�7�t��"O>�����Y�ݺD�^l"O~��ۺ���{�M͒y�>���"O\��KK1X"`b ,�<� �"O�8�S��?Df �1�90oN<�!"O2�2a��9�A��1@p �*D"O�p�� @r ���U���!D"O�(��"ѱGXX r)-:	�T�"O��
��RF�LT���j�2ѣ�"O�0sQ�˳Vx��3�LK1W�Ʊ�P"OFB��bS`ٸ#A�L�<!1�"O`	`B��;!�(�� �]T� ��"O��i�Y��bd��1DP0,;�"ODT0�FK8N�L!� Jݥ*��[�"O\d�ʬP��'H2c����"Or����ʛ��݃R�߯X8| j1"O,�;� �}K��p�FQ�~'�H��"O"m���+w��H��2 �jb"OZ=!�j�Tm�f Jh���s"O��Si��=������Nv��F"O��ki��?�QR�*U��E�"O^�rf�C3De0F��
��ٓow!�$"'�l����,b�4h��@I6A�!�]�K�	��g�
 8tE�)Z{!�D=� ���I�-�
��e\�E�!�D��W}����a_6_L�@��D�+!�$�2AF��D>e�U"wB��!�͜@ ��(��.+.�`v@� !򤎖&�xІm	K��Hy�V5f!��Z1S�萃��J��}( -��!�D�	��!��'�,U�����[�!�>]\�;.��Ih�=C�(Y�Nu!�$P�&n6d�G�.MP����(N)of!�dO.q�
;�ߟxFPa�c�3e{!�݁[m�������*�h��T�[r!�D�H����p��e	�0��Nl!�d��B:��z�ϑ�M�$��1c!��O�3w�l�F�M�7l�XKS� �!��](>��Mt���Qj�0B��^)9�!�d\��MQ�)\L(��$�O!��q�@S�K�}7��3�� ]!��T5#�~ ��%ַ[�����_"G!�d��v$E���R��r���W!���"ߴCô����]8vڀ��ȓ.�Q�덉t��Ї��1-b���;&�	�פY)e��pGO��z4����')�0��N�g�����Y+X�u�ȓ#� �[�Ҏ��'��&[�L��(X��y L�A���HGB�f�Ȅȓt&\:E�"$A��@��]�����}R���A��?���e��f�&l�ȓ%u��`@�ʈN��%�vA($#d�ȓo"� �9D�0�G#F�4ر�ȓJ�x�SmO����Kg�A�:���@E���i���F^�4X���q�l���K<��{�m�1J�����r5�Â�'�J���nG������G�C�S�^���i�$8����)E�p{���cd�}Âl��g�ƍ��~��9Bn�)wG�����7Q���h�"��Eߌ�,1a3o^�;<���z�H�P�N��`��D���M��-?�Q��aJ�ȝ�ቍZ���ȓJf�ɸQ�Sǚ�r1}�����S�? �y���՗dN�=;�+��"�!�e"O�����K{~����I�YFTZ�"OJ�
3��!I�8$Y������
�"Oحa�i��<�0�J�S	 ��"O$��B�7�z��c�&L��S�"OV`3L��vaz�0�	-)ʢ@k�"O�<���C=���Zc��!��й"O�xbl*a
��� �>Mh�"O^�S�eZ.p�h��}	��E"O`��� e�݁2�@%%b�Ix"O��`���FOL@�V<Y���"O��
ˆyF��ѷ �)Lפ���"Olh�o45�̑s�JҐs���"OT�j4�P�H�˜4QR�B�"O � ��E6\�@ݺ��-f.�a�e"O�a�J�?Swn-6
S�&)0�"O�Q9�Y9o�#P�ґH ��"Of�a�.ҦxD<��Ԕn��X�"O4`r�$���`	����'V8�]K"Ox9D���32��"q��<{�N��2"O��"�m�X��%�^c`�Ʒ�yR&�'	�l�Xgӏ1L�#�C���y�o�0X��5�&)���%����:�y�mC7'��C��_�����&�y�F��(�RY*��V�P]S��y���B�,8êHp:�(� ȡ�y��	P��t���]1B�n����y��Lz���Rc(��U<�yRf��]Ռ�J�nƴHp�=�����yB��5����.�X�nu8��U��yb�f�X�xV��|L䕹��A �y2�O'�M�ޤr���aꝊ�yb��"P��{tbO�2��XjVB�y�)B�T�c���/E>��ݖ�y�ʖ(wF��h��'�=�!Ǟ�y�`�q�9q���-� 
!H�<�y�lP-F����m��	$�S�g��y�+֘	 �4�GJV�ܱ(��y�Θ�S��Q�.I  /V��y�-��>5���9�����Ƅ��y2��<c�tBV�Ј=��q3E�Ҽ�y�)�z�^}1��G4�N�JT"�.�yaC$
�j��0�33G%S�0�y"�T}d�͋>\\��"֢�yB��5F"ų�`> M~̊�	!�y��V���dTn�8̘��#�y���QP��2BJc��Xdl��y���"S�q��E�C�ʙ�#(X�y"-�_��}b` S{|���X?�y�E5� ��	&N讈�v���y*�M��DX�o�AE�e �/�y�E�J	9��&ݨ�b�(�y�C9V�@m "��	*<\ԁU2�y޼'�qyF��Y<9S�R��yb�ΟlR�]1�Lq��K2���yb�Egm�(���\ VD��1�ٝ�y��6EVfl����&����Y��y��?����$�fn��Qk��y"EP�H`x�:��؀{��<iQCC�yi�+�(�2ĊC�s8ء`�G�4�yRψ�.�(Q���\�g�p�ʕK���yBnU�#.�Q���ūW�*��E��y͞"p�
��i Z�=��(�y��5S��v�̗G���q4b���y
� (d��d�-^x�Ő�j�:G�����"O���`M�b���ʠ� �yuP騴"O����a`�	C�\���"O��a�B1>l<���ܙcv�� �"O�AY�C(����H�|9L�z!"O�̊��9nh��RV>{n�[R"O!:Tc[solx��5�@�X�"Op5y.E�:4��o��R��0ȃ"O��d��9��ǆ�Ev�q�"Ob�8 "Ʋ<t�z�g�c��L��"O   ����I"ڴ�ԦJ�gЙy�"O�U��'�8P�t�aE���l�i'"O��2T!0^�r�q��h���"O,��n@
a n8b�Ɠc򀐐q"O ����R ��G��34�0c�"O�̓�CA8a���ȣ �+���V"OHEj2��
%l�Ȁ�� 8� ���"Oj��Cf�+wĎ�  L3d��@u"OZ�#�d� 	���U8:ap}q�"OZ4�k�0?4)���#N~��q"OB��1M׭s#8�qƠ�Y��A&"O�İAT�D44�Jc�[
�ܨ�0"O�P��mC
\�V��a��u�V��"O�(׌�%��Z`�.I̼�JE"O<�
��~�
As$	
8F����"O�9)a�ƩKID ���پG9�d�!"O���C�H�Q$�@i2�	��"O
Hd.N4[1�8��,��!V@�"O��8���p��s����usz��"O�X���8e�Б�o�	D8F�K$"O��� �W=r6�� a�0=ҽС"O��HF@X8Q���&{-���"O��Xe�ի*�@dSԄ/J�p"O��Ye	�p�B�3uDܓJq����"OPYvH�9c8�ܪ%B3k�L 1"O�H�O�d*�q��D¶n�a"O�H���N��2�dЧ:�d�"�"O�	��$��-�TX��DY�b2��"O���F�y��9��׌o�\�00"O,�����0���B�ۈ0���{U"O�d�����4����N$����"O�R��P��p���]8��7"O�}�$�F�$p~�a��#i�YA7"O�!��j� KPYTJ 4 ���!"OXa�.J8r`P!iّ/C
��V"O�x��
���Ia(ɡL�=x"O4��&4BzGh�RD��6"O�dD�
2Xb(��-�)ta��"O*�a�nx\��Bm23-��"O�Lj���� �	a2暬C�`�"Ob�c��ұP�J��q�ƨV&�Y�D"O�-�o? q��?2H�Z�"O�䋧��6Ʉ�I��@L~��@"O���*DK*�q�`֨^i �W"O��'��o�6��A�<mg2Q
T"OtP�!-[&R�踈��[�C�Ƅ��"O�i��KU�<h��Qp�;,�Rx��"O1cag �z�~�#�,�9x���4"O�� dDV?$��&�]|���"O�D��
�<a�䢠B��6R~|�"O ̫׆F�RP25�ک�F)�G"O@p��2�8��wc	6u䤂c"O,���I�'J��$b��J�mdl�0"O4%��`����k��w�x��"O� @y��Ђ#��X �K�.� ��"O��c�D����!��/��I'"O�%���B�[��8�N�(�E�g"O���r��6e:칃��4>�L*a"O�Q;��	 s�Dx���MM3Jx�%"O<ի3��!f҄xW<=(<�Ҧ"OT��d� &A�Q���X�7Ф"O�HAtNԊ?Q�� %N%Nz Z�"Oޥ8��/:�����ޮ+5�Y�"O�-`֎Q�����F՞(��-�!"O�c�I�$w�`H�#�A�N��hh@"Oz<J��Ճ�m@����e��h�"O���UA�E��G��X�h"�"O�=��@ޗ3�Q�늬	��K�"O�g�Ї*�e��)c}���#"O0��� �o¸	�%ȇ�2E(͠�"OP5
2苊"4�����[�Z%r�"OTM�e�\�u$�1�g`͝��9�"O��x�'&�$#�¯����g"OB�#�-F�J�i�nY�d��ᙅ"O�Y��m�K*�!��0d��P8�"O�p��V/GMP�"�ތZ"O���ծ�<�(G
���`0R"Oި�% J�v�҅b�,�o��u��"O�����ўK�$P��[�C��ݚ�"OP��&�scb� �+q��U"O��� �ƘgD�J��$��b"O����L4@�2����Wuz0�W"O�(�r��>w�V��B���Ao�8��"O�1	�f5�l��ċ&P���"Oz[�!��s�t`c!)[ް)��"O��bsŌ�h���胬��є"O ���q�;���	'�h�&"O`8r�D��G��b%o:!��I!�"O���π.)�0�#�-'9���p�"OL��  �?� !�P�9�9"O�1A���?}���Ѭ˗!�L j�"O�I��-�� ɛ�k/�j2�"O�|��[�G"
��R����"Oy�bF�P՞�U�PUI�V"O�\ ��A(K�2Xpc�f�XK�"Oִbe�>o�4M�$�֐?� �f"ONp3�@1g�~�KE腼���1!�N�	V=�`Ɩ�H� eXc+��Y#!�Ħ�(pG@}Bl �T'[e!���,{��	�a�qs�J���Z!�$۞g��@ۂF�@��I8T&#@!�d�#F:B��a�w��k&P�r[!�$�25"��'F��zi��ER�!��<���	6�
� rt�E+y�!��̥co��A�i+G�k���2�!��ܬX�8
��ɜE<||ꑈ�[U�'�D��I�t�(E �MU.P��cʱ��B��Lp�5+�4Z~�s&��;	��'�ў�?)�2�M�+����,�8nH �R��:D�����I7v� p"K[5c��`fC�>��)ҧ2�h'�(]�@��9^�����m�~��-	� }�Yc�HY����%�h��I�m{���hB0x�.ٙ�ֆ����D#ғ[5~�9�GA3Hw�d�P+?`D�Ɠ�6�#��iB�뇫_�LH��	�'E�q+�1{��
$��K���(�'�P���ɇ`n���"@�6ي�'�pպ�
$P�v�Z�Z�%�f���� >��� Q�$�&Mj��^�O-(�B�"O4��`i�.�V��Jίk�,PE"O�9@� ׏p2����i�{�А�"O�%���Ǡ~�ҩ��G���>��{"�I�4Hdh��>'{؁�Hͯ�*݆�	I�I�jЌ(��7L�m����zF��hO�>�*�mG�1�h�.2�R���b3D�(�f�Z6%���*�9p��q(=D�\ȓ'_X���C"T�M �z�7�O�9��|7�����Ea�AJ�)�ql����ēdF�#>�'�H�jˏ`St�q��U,~v�,Ӊy\����[��<��kH�&�<h���[]}(fę+�0<Y��ʽ�$��'�#@��ҥ��-IvB6�7������X�'���ꇋH4�"`
�lJ�Pl0�'� ��բşoy}��mΟq�n��
�'
v���"S��.Ukb��2pE�	j�{��)�	@��w�˴:�`<(%l�<F��a�:����w��v+��1� �!�'��'C��r���O
ͫ���V:,�����'�jXC���;6��իGC^�cNv�X��$���Й���H���hr����-�Ş_�����<-�])S̬8O.��Y��(�'�]��n�6�\"�>�E~��d.B�o�Pp�n]��P�H$�[�<���C�7��q���;=j�PdFQ�'1� �O�T�rf�fm"�ڻ}�Ѐ��'Y�M���A�L4Cm�|J�)�A�iZ�"~Γ��ɓ���Y`<� �J�d�6Y�?���~R1�\�UD9�ڄUSt9�ÁX}R�'��5S����jp�ȅ$� � 
�'I�����_*�z��>O
�+�'~49�6�ӂ�H�Y�BZ����1�Y��%�2&抺D^M��"O����&�*o7"\�$e֐��p:q�i��)�禵R��:4#2�SR�˅j�~`臃'D��8$�E�@f��V̈�hlBR��>ɳOc��=�}���V�d�`�)؏Q[~�0U'S8��IZ}���"5�\�@�B�����(��yL�R��cU���|�j�OL.�y2����њt��
B�4᷀��p>iN<�2�A;EĪ�:�'� f��+��Y�<a"EX�k"��q���}J�ysV#�j�'@ўʧ���r#λ9J\��?�H���'铮?E��'D���K�T���bmRNdFP
�'I|D�Ũ�,�4ZW��A�f���D&,O�,ӕ�
 {���Mo�!���'��'���M_4n�|r`aD�}Dj��*/$��)�DJ�&�̍�ć���*q�`.*y��<�O�@�
+���bg+�I�X�9�'Z�y��hZ�cj^��ٵ,\����y��)�S0��ɳ��9�p�
᫇� ��"<	�>�S��i�Ǌ��_6k:M�r"�!!��B䉷]<��ԄV�� ���@B�by[������ۈ���Z5K�,�xM��%o��}Q���Jyb���y�6�4	Z1Pu���t�ʰD���y��u��$Ţ-��xp���X�RXꔄ�{������Ex��	�21(�3%��>�:D{���,�1O���,��'�'3B"gCK'��-�4g�q�'Ŗ�We<���!�oվ'�����'����C�����'$*��4�Px���29v-��MY`&���b\�M[���'��|Rc$�7D���G�"��	b�'"���B3(��c'��|}z�'o�S(�%J��u*���t��O��=E�� ���1�]�=~�dۡ|bMpr"On��㎝�l��������R���"O�ERa���Ī��F�5�*t�`�Zj�8�'�إ!��V���x���f*B�J�'!ў�I�@M�"N�r�EI\@���*�d�7��'q�d��N{�	�e��<�4|c%�&�O07��<��Gα��=)E�
�y�p�hIC?)�Ox��N?Ɍ��'�X�P��+��&F�$x��،��|�Ԣ~R�/�`�X�gɚ�g�n����N[�<)�,*J,�jvQpvԸ"�o��P��I�<�.E�6����#��<I�d"P�h�������:'�"ŉ����Y�+
��!�dY5)#jy���)n����D��<Yy�\�W�)
B������� �M���H�O	a�<�%G�n^�jpC�00B�1���s�<y@���}��`aLH�M�T8d��f�<nȘk@m����&'����u��|�<��CO�>������a2B��DǔA�<iP#�)xP�\4��c4�a�V�<��
?/�e��G�9OY�)��HU�<95Nܷ! H��DH��]�A��jR�<���_�xۂ�ƳQ�<����I�<9�-+op!�e�
p�𻐎@�<a�jW�@�j|a�O,	蔘k��x�<�F�E ��Q���#����r�<��B�H��<�A��#$քQ:"�o�<�S��'[P�s��æDq3��(D�\)��$<d� �/��"�%D���M֕8��#=`��AA(D�XQ*C�[�����O%Mh�9�D`$D�|�q�95v�#�B[�k��6D�b�ɓ�A�Jm���2��8�K7D����ʷY&�Y1*	���[&h3D��mM�N���1OF�7�����3D���E����R5�qq8P�F0D�`�L�*Έ�6c@"C�,仃(#D���BG�^�y������{�mn����*N�9��N(�u�T�^���'������n��\�	�����'e�9y�%Ԍ,�(Xl��Q�ݴ��'�l�)�3}���x=���m=f��2W~؟<�����c�Y�i��d)a��q͘�s�OZ�i��;X��@O��C"�x[��'��O�p�ƍ�/s*p ʲ��$6F�;�"O��*��T`h8���!�v��A�"O"�i�mTu�-���T�m�Ι{v"Olm�A�5r��tã�Ŋ5H��"OvY��F'1V��E�T8/���i��'�Ě9�| �ʌb5�}�#'�N!��N�~Ò` 	�% ((�p윴A=!��3=� ( F�N��J��#!��?p.�:V/���Ѡ(O�!!�$(:2`;ӌ���hXrR��T�!��:�,���7k���%�cH!�O?�zM#fM+.���I�k0!�/�,i��Ǻ��d!�C�:)!�P8k�EYT��=��L�$��X!!�E7H��q�G�-%�������'!�D�#9�[��ܠK4X��OE��!�dɣsP��A*Z�oT��aϸr�!�R$6"��cd�]&�=2��C?���_3������ ~5��:p%���y�Ð�k�F��o��s="-y�Nȇ�y"��"ܖ8�aɁ]���ֆE��y
� ��fb�0i|N!�dԮ`�5SE"O*����y�b�r���8��l��"O�LЩ{�ݒ7
@�h�8s"O~`8�h�2F��"%"����E�b"O��H%Dɬ5Y`�Kp�I/a�$�Z�"O���IK�n`�AS4O��~ZE� "O>�3� @�zE�V���G����A"O�hs�o^'�D��Ԭ��B�&!�&"O̼8��
�����d�<��"O�����S�+/�4X�-G3n�U�t"O�Da��2c�"�P78�f��"O<݀�Ҁ(�|-CL�}5(T�%"OdÁ��4��F��<b�d�S0"O*��Ui�*��8c2�1����"OXM�AE�wp
���g8���!�"Odl�t��1"
�ؔL��h��\E"OL��g�E�F�i �ղt�����"O�\ر��7l2�lc��>� �5"O��¶"��c�*���Ź.��)�"OjH
�S�rՔ��5řn-��"O��K����� �3d\�Q*��y�"OX�S�Gׂ����6�Ǆ���!S"O89��,)3N�m�����"O�г�N[/=���R�F��jJ`"O���iM�Q��m�2�Ni�Bm��"O>�Ad#R�V�p�pbWW6D�ٱB�C9<���' �`��b$\�5nc;�z�rT�!D�@夑�G�B,�2%��,�$@��-:D�к`,Ŧ_���'E��0�`5,D�`�._#!Ϯ�w���܋��*D��歛�FW��w��q��Dy%*O&a������k3�ż _f���"O��&�ZX
���Z0�2"O��!`�B�P���F�Q2w�$y#�"O2<�g疢efzx�d4V�Zy��"O҉��ˁ�;r	*$ܝ��"O�S(#-�H��O�6�@4�"OR���@=�.�<x�JX�"O��Rb� Q,�m��#5]F.�4"O6�)$%�q�d ���ߎ/>|�"ON��Tg�L�Zr��RPaȑ"O�3W⊭rfE@F��9�,u�"O��;rNܺI�\L�b^�f��p�"O
�6�ėB� ����s���3�"Ope`��%��H�1)Ҥ� ��D"OH�)��K�P��|�ዕ�v�8H��"O`�X�K N���hP(0Ūp��'� ���$�9.�ɧ��z	v`Q�SP�O�|�T�d�;D���R�2|H��P�є5�J����>�cJ����At"$<O�$�4!QHT��ic����'Q��!�ό�*N(Y���t���+Ұw8T1�P�*!�D�/^��EJ��BP��8�Q�X�3L*J��%ʒR�'}�\��gP9 �t����� K*��ȓS��J�{G4=��I�:�L�:ş�Q4XѷL��)�矜K�nK�iN����،pD�x M3D���s��?i�59?h�ҥB77��	4Y�8����Ǔ+����I%FNH��ែ=^�Q���h������XֺAc�	�\~%ffK�^e��yc
�b*h�B��7$��#KV2��tӂb!%r,�0�h"�"�*�K��0��dÊ�de\y�DD��	������y"LA�H�|j3�	@��dإ�Ֆ ��4&5���(T�<E��8��*�ǒ<'p�|��a�d�0%�ȓ3]� �!f\�J�m�� ��U�\i�'��E���=����!��pGF �$5)Cʆ�KT����JP5 2�*� ���T��(��)5
̟A/&�h��'��bP*�S�a|A� &(�g��[_����T#��=q@k˹=e^�J'�Oy��,#f��I����r"O<8S4jU�,� e\�l�ބj����6FiL���!#S��"}ҐK�:�"�yv)M�m\�P�7i�b��Қ/ټh�O2���հn��e)T@�9���c�"L�H%�f(ٔFL�'�8IG�,O�`Q"n ��e@�G�g|P�6g����Y�2��.�3�� H�z���}`���&b�.\��M��l<2����.�p<�ҵj�� ȸH�|U��	�q�<�Ѧ�)}�������""��z�M�3h�6���x=���)5掑CUΑ>u�џ�hÒ*���{&��y��ۮyR�����ҥcWh��̸'�ح{t�@��b��铧|��|�B선&�J�X�ܘ+��ʓ���J���ui�D�
ç|�p]#��)�l�I���7NV7�p	��Z�`xS�<1��D'cĚP��+G�n?��!�m�&@|�'���p�fI4"?�ϸ'� s��&V�0#C��^�D���n��%��q�E��0h�<C�V_�@�����#�p�sAH()���Â�� `%��*���<�����D�xDց�?�E(�	w�����	��6�t��T��A�]#:AZ&�V�:%�ݺ�f�%]��$�5�?�F͖�=��@�R�0r�F���<���4f�+���m�OX4T 1�ٕ<N�=�'.؁��t(楃���E��Z����O��(��| �'2td��e�$�P��Үj5Jm�'LM�C�4Tɒh �.g��i���%;�e5l�Sdj�Z�Oڗ\H]F}��Ц0T�ҟ%Y�Ȕ&
�O�LP�jS!��Ē&SŨT���V�
e����"�(Ā`��B�EAҎD{�8��"�Oti�t�1���G�[g�������H��� ��O�,sU,�/+�,y��'�ּ�6�/����LL4D��CV_N�<�DG\}Ӵ�k%%Ȳ6��|(��Ox�홗��WV�$c�'�d��qw�U�vNU�����#@6w�4cC�y�t܄�	�dj���	BGTz�jU��YD�Jw�$t�1qeᆨS�.���=lO����νu1��0�*N-��D�b����9���G���yb���;���c�ʬx?���*Ѥ���@إ��.!G�4q�' $i8'_�ItZ=���� �$�v�$|��d�On�����<�����{ޭZ�ؾRT�4���\�,p\#l6D���&W�.^����^�\��� ym|�Ƀ9��u�'���/W�$Ex2�ؘUJ��
�\?\�Z89"��ϰ=�ǋW	"-Td�)�OVu�׌B�� �0D�öU
�)2v"ON5gS�*���C�8

ɢ��@��`����h���2�� 8a�����}����"O8q���$:*&]/)�I	G��=_�}pP�OxAq����yჅ��?:6f�/(��T5��-j�E�Q1.�kd��5aĄx�"O	b���N��Z�%�&���;Ph�!4ˢ�ؔ �O�`
����O��R�O�� �wc��h�#
A����!��p�Ĉh�'�f�CŖ.ij� �����P e�ր8Vf����,�҉A�NE#R!b�3%Vo�'��`���"$����Y,w`��;	�%����3�X.th��k��
}9�ف���x�"���?M|Pу����i2�Olt[�˘�Z�)ӷ�C[T`I��|��WLP�G�#���3�E]3xW"t���V��oԾJ�R2���%��%*�g
��y�oӘG	��Xf��=�jɹQ�ʦ2�.�A4�]�cl��#pL�?�lr�/3�SR"�ͻo�c�H��NWLm��Q�w_���Ɠa��|y��5\Hأe=���tn��x�e�>\<N���,L��T0A)�We�,yE�!��u�Ƭ�ƸЅ�I#��]�f�U̬�15&O�F����C>6�jRDR=6<�I���D�(�C��'\̔���L�F<m�C���}��4�O>�c+~��,�%��Y��l1@dS�:�f���H�~�YYF��2�&����7u�<��ȟ�#y
���ݒ,�@�G�_�K��a��M�-�ͥz�������F�p�X�]_d�r��u��8��L�?R�B��/��5)a��J��xB�ٕh�H�GG`��.Kx8)��ʍ4@ ݳ�M����O�Șg�^0G�5� F̼StL]97�'��v�5�F��'����Gi��`���L���Y���'� ����86�|42C����fΧW.�'9��c�̟J6�T���G�f����[9`9���O9���+ r��i��O5b�
���'餩aA�Px�f��5]Z��2��5�)� Wj��d����>��O������<�B�'=�иB���i`�@��BHM(<�&"�EVb�sХS>$�h�q�#�L�X��嗽X>�k�n�t;��tDCZz#>���0���5����6�A�	S8�ȸ��W&C8f󔇅'PFlP��� ����n�����B ��#~~L��#���BŁ1�'tzVb	/R/Nh��Es�H���F�߹3�� 0��C�F�R�5��
k���+��?E �+W}6	����;�Z�q�M!D����Z� �ȕ��(@?^5�)��o*�E0���Y��PEP� �b?}A�����y"C�8��H��L߁ ��T)�����xGT�j#�y��k×�$�1�O^�L��V�n�"`)A�ff�Hٵ�
h$Q���fb��y�xy�Ҧ 펽��&R,!�򰊇��Q�'��k6���M����c*��W�`������s'�kĚ�Yu�V}{"�<ٗ��
��S/,}�.�)N4�����.j�扊�ۈ��'�N�X3��s&Bm��_�9�rY#%��tbN���0R���4����$�Tfz\xblR%l|���)�'�$U*��.nѸ���'\��*HӤ rɑ��v��X��<I�HO�>]\�£%D� I �lS�`��\�'R��AͰH��ϸ'Tj����<0޽�3���-�F��{����cC]�;�4�A���Z�d���S�Щ��h�R��D��M��fY<;	�a�,�Z~�4
��½�~����e���y��3 �:OL��O����g�X�t���<��.P������\�8s��B �Sg�Z
�|�T�=���P���#l	�L1�Ác��5�'��9��EA��!���O]fH1c흿?��hg��|E+O��փI��=�` ��+�t �/��U!��JP� З',^�x�)D���M3�łS��i  ����|9�`�V�:4&�sqdB�v#b��*�r�br���e�d*���"�R�B5N�%��0sVn�<AUK�d���z�����c?)8W��}5���-^�^� V�7O���*�`�RN�\Z' (\D�3 ���q&,%t���`�>��eP�'�f#}�'N�l��B�1h ��k��a>�d�N��PB-W$*�x%��?����AOA��7D� �2$Bc�<0h������� `#W�& B���Ғ�a�`˃ �`q� �(�z�Ĉ,]�4��) p\e�ˌ7�>L�QGK?��t���۾SE�Ȅ��|F�	��@8�pAhB@Ԩ,h���=1�7���cr�:`Υ��K"�S�El	���5|_NL	R��	p8B�	*
�@m�a�*s:��LD�����P*U�=��GÑm�@��j?�'��V^��!5@[?+ �းO�!�[9V�tS0��+P�`��b�d�1�L�9<�b�oǟ+�]`6�;�����鐏<�@���HO�:B��	X�������ʞ�W���hf��8f5D��!�3K^]#��dr΍����<j�K�f<9>�����o/�c���Agєk%��I1cG>fFݻ���i�ӕ2i�a0geƬ.� ��7�C�l&B�I&L��y�vÒ�|��	���M"Pz�y�4�j96	��\!-��$�'>�'�򄝫aNZ�[��	�j��$�2�!�$G4a���5`N�"���B��y�r�aC捞X	���dJ�
O �'�f�5��͡m���*�툅)IL\��6Mx|���C!-��x�O�p�4���B��9��A���r�0����y�Ht
Es(����#�"E���X����[y�����S.��[����&Vvh�ժ��	l��[�!��`�!�$��">vm�CLC${&��Q�Ѫ�ڜ�c֤:�$X�7�� �*@�<AR�I �x�a�!|@zg��i�<qDJW�BY��X�"і�̕�MQ�*� -��3�@y����I	}\�H�؍�Ш��K���$ޕ�T��!I�!��h����+.:5�6�{?�l���Ә}�C�	�T)ԙڰ�h�@Yp#��_����Z�+=�Z����ѱ��pP	�4o��u�ǤߛE�)S"O, "!���q�"#��W�T���B p�%'n�!30�S��?I *A�FR� �F,��dL��	0��V�<i��B)x�2P����-���8ӧNyR	_7W�L��	��� �`��n��(4
��4�C�I'
]����瘿0��w�ƞ\g�C�	�h���xB�Z:M:����X.v�C�	�@<	G�� �B\B����FC�I,)ej���k�}N$�O�z*C�	|�tC �Pܵ�WM�	��B�	K�i	��0��	PnR�9�B�ɲ%� 6i� <Ebiӣ*P�7e\B�	\Mr� �"�/L\���u�S8G�XB�I,n��jS&�h�����/�hC�ɮ(�d�bT�FRT�z�F�'Mf8C�)� ��z����,��LJ �	.C�53"OD�s�<?�\(�����mD�E�"O��_-#5|��9�q "O,�AƁR�!h�ъ���j#p��"O�:� ?N\>�!R�;{�"O���	]��t�s��A���"Ox�K`��E�4)b#��0B����"Or5��A�9�L�S,�/	ĵ�"O�Q�QnAv���F��E�xH�U"OX���,W�J����@��4�( '"OVqK�<>�4{R�¸0ҍ�@"O �92�s�|��Q�s(�t�"O�<ah^&.]�T�ͤ;&~,��"OL��#NҨ�Х��Q{<8��"O�� �	(�`-���V�-���H1"O��4�;���a�18��!(�"O�aꂹ*ipwmE������m�s�<��D;@l"U�p�Bq��MWj�<�a.(X���4�t��Sí�\�<y�JU!g��CSL A��A��AZ�<颪J%{���= 8ڀ��U�<��g]u��9g���G��<C��P�<��e�0[��`lC�?�t�R�͔N�<IV#МJc�U��Ό(,�(xu*F�<���#5�M���\�k�:��-|�<A�B��3���*���))�ƨ���D�<�Q�S}0�Mr� ���zF$�F�<�J�#:�HY�$� �3�+T��2`	�p�l�2Á�bw&����?D��0��P�`9�PQ��#] $=D��؁ ��u�rx��)�&b����=D�$�&�ĸ*(���`O
(�lk�F$D���f�\�k����J8��I�U�6D�p�c�s�Ψ���կX;�9�8D����L�DN���/�^fj4D�(͒-{��42���$��ys2D��ҕ商n�42��:��G�2D�L�VD�;%pɹd�Ѳ[����2D���+͘/�Ψ��@Q8��7�0D��rfn�?�*���)�!?T�"e*D�y�ˡ6Ox��_VB�!E/?D�X1�M�pZ`�uX�8�` D��bF�=	l�� ��Y0$|	#!D��@��ͬi�)�cA9�� K3D�8n'���艱+G9,	�lcEO*D����Ӫ:���@�Ѽ]����%?D�谰�Qአo����y���?D����O�&]�g&��.�����=D�l;D�¬K�B ��$T.u�9ic�)D� �W$|C�
2��,��=��%D��$�.W
�@�EG���Fi�?���K�:T`�I>E��H.H���eM9y(�!S��� �!�ĔP�X��ڨ,s� �o3y���W�Lq�3�	y��y�k��U�����3y���F�ۙ�p>����m`��b�I��J!�c~���t��Y�����'��1K1k�$$����!���^ÄT���H�Y���+�&'��c?���^�T&�MXR�E�[�Dm��b#D���`�%M��ca�0v�z&�� H(8�:��s/O?������B�R<@�<��
�!�$U,	���#��4Z �d�&�"Si��Н:d�8լQ��'*�7(������rW4�P2��b8�T�`Ȼh�L�Y�'\�BL"G�/q^�:��.~�Dy���ԑ)Q&X���� �'�HpGy"�6���y�&ٜ�����@�2�؈Y%@��V4X��"O� ����� Ұ����ڽ=$$���k��d9R�*\
�ٗ���B�
�F����S�r���������y���66r���2<x���g����;���s�h����<�P��� �����[lI{��gx�Lk���'
�ca��d�R��oP�V>*��4)�ݟl[k�*
���	!Z��Q���2&:: �#� 4����d�s�I(�Ґ�?Q��Ү"��S�T�,���+$�v�<agE1y`�+�L�!M�`��ɖTܓW�����ʊ;-��Ë�iZ�#��݈���9b�4�8��J�c�s�a*Q���S��k$Ё�!˯A�hcf��0`F��B�
Ƞ�:P��9e�<��
�9��9��42 ��m�nr��'i`�i훍��Ϙ'�.2w��NY<X�B��/&!Z��@��p��TE'+qj���)��͠�Ʉ\���K�G�N@d���� �i�B��5,+�u�v�����,GĈ�4��!s�ɍ4�2@1i�	>�^�GBL<"=�� D�{%�S�6}̽��-^�l��i7��2\ߔ㞼3�"�i�J��N�u�O��a��a�&����"͒�|��#(O��Vc�7M.��3p� �̔�֠ǁv+�m��^=�{n�@;p�A��2ʓ ,�|�'��=x�IݢBo���SOÌ-�� �����d�9�8@�"#���JƦ�`r�����@�6>����Ұj$���D07�Q� c3��?�
�+��ӳ_�Y���
�y��ѕd�($��&Z�T�F~B@͚-��0�a��2�˖63]t��	
-}�D1#�O7�I)P���%h�.Z��T��b�&-���͟�y�����͚t� �]�F����d_�Zxx�f?�0f0Id�^0	_�iY�� 56��]�p��G�����\v[ LSCi�d�O��I�!E��TCF�K�.�T*:&a01�ȓ�΅��@��N+Ľ9ztk��h�N�"���
"W�͋s 64����6�	%`���{*[3���
@1�"<! b�K�P���G�A;�D�
�|j��Ǩ���D����B#~�@�����8��?�!$��UlL��%1hT����F�Lp���t?�C��.�p2$�+��O�.�NFN�1BE��6( T`.9|!�2�^�H���oq���q�\�E�ޠI��Db����6�j��p����LS��٧m&�O2�r�Ɲ6=�p'k�/2�"����'�l��چsR�l���^� ]b�J!J�(���
�0᮸����'��<�J�ް=AӁҭYt^}H��E�~S$H��MUL�W�D3Ճ̅I�b牎��Q�P
7V4�p�;L�d9+Q��f�P�T�V����'�t��iN28̸!G�ԀL������,��8k��Ol��L֯D?v���tKw��vMZ�~����.)�a�F4D�P�F��;�� 9�%��I���Gc�%@n\����f_H��'��̓
}��Exr���hj��f���-��g��Ӱ=��cS�X�c4��O|  $֊N2\��!6��q�"O��C���Z6y����;-::����L���1����h���R�� Mi
- �'C�	ʴ�"OQq F�(GF����؉1�^��� �gNX�b�OL��ע_צYa ��?����X�0���0��E�d
�m��(BB,8���P5"O��x��'h��4�#A�FO�lhbh��bm���O�IH���&�����'i��<��Oh2$�ws�l�t��-SHd�1O��EP�'�f4Q�`�^�hs��8]g�$�$��u��0��K�T���e�Oub a��N�'� ęWf�5(}:9Ag%�87�*U��)y6�e�:4�>}���@�xvE`�3?��]�H�!H�$�Wsj��sN>�O܍�El.{��:�/��F�I��|�Q�J�yؓ�ܛ[Ȣ��'+@�F�
�(�D�ti��q)F �@@ӊaaLP���ϭ�y���(-���(a��V�����)ġ�"�]���eXQ�U�1|���=���&���wg
u�e��-l���G��x��	�'�����T(<]t �$�I�O��)��8�X����M���Ҵ�ޙg ����/Uk�'��\�k�O�hѢ�'u�)yϓN�d���%}�)T�̈́1>��e��}���K��N�ؠ��]�H@�w�>�ON��0�װ��Y��@6Md��0��|� [7Nc�� �-���v��ޔ	�}���H�&�&���B���w~a����y�ľ|�>t2e
�lCtp`@6JyJ��7H�Q�$��&G�� `����� a�Eλqx�G�נ:a��R�ڵE���<� :��?�$9;��_��M�^��`$K��]�����ʉ�e�"UC�G��H"�R�8/|;p#Ѩ3���#-O� p�A�A�����O�Q�s�ٳgDX���$&n�eK��=�)[f�%�O��⃊>z����w�H��>�s��%��-�k��= Dt@�現?%nlz�.=jL�`>9�F�'4����V�<� �x��_��~�	s��)k�ᘡnI������LG�2����`��q�JM3���y�/J#82FCR.�r$ h��Px2�G�z���S�O�"D�T�,O<ƙr�V9=*:��肵L�"Ԣ�*B�b�G|2�T|�h�� `eؙ���E4�p<)bU�+��Q7*V��eb��;�M���;K�T��ω0K������X6*�,���_�e� xjB�8�T���D�\��Zs
�8'�	u���3�IG&��Շ�sPT�'Y!pA�$D�;ٶ��v(ʹ
��Ɇ�x���`$&d✌`%�N�����g�bGFP:�	R���k�Xh�;�J$
6:O�x�A�ӌq<h���_�D���&O�x	t�Ѹ�����G�)��[$	�C��+�Oѝh7f�1b[<F��q$1�A�����̭`��
1`�C�`1nXd���ĉ7)Vh����dάA���K�6X`�� �+��2d�L(����-�E�'�6LH�A@*)�쬦O�(Xpo �8�I�G��?_4������,�j�	`�Ax����=^���<�.�8Fd��R"܇.�|�r$X�t�UG�s��¥��`>Q�#͜�.�(�X��C�y#$5�q�=��Y��+�g*:�͓�ң|�',�%�G�E�wx9Pi�ts(8�FZ��@�^k���@�:��D��d����ݾ<��(Z�-�n�YF��*����C��4�џ�: $2,<P�S�O�0�&�1�۹���D;0���F~"��k�Ľ`�O \�e e���c3�\�p{`{���3���3o�w����O��qР�J�@��`Cʑ�3
|�1�b/0�9G���ŒWĵiu P.�P�Jd/��䕀C[�X"��?om���0�Y*��̆B H�A`_��!��G"�HJ�G9�`�һ=n$��A�"�򤂸I���1�/��$��A)Č�FDF�p�ƭ8o]CB�2dܧB.(yʒE�3�8!zt�W�z�q��mR&/^HL �'�*��� �5ɈE�L�yu\l	Ó���`���:b��'˜ii�͖E�JP�թ�0@��T��'�$TtK��gi5Q�	ͿmU�O�,z�
��~ٮ�'��?��ώiVH�ae!7ql-lRS�<1r�S8~��j5�D".߶5���W�<�� 7Ez�ȱƣN�3C�5)G�R�<�'�M'e�0ɡ�K���0�E�<�)�aJ|�H��C/��� k�<Q�� Rrb ��oXH�Hy��b�<��ŗ�4|"�҄��`�M���PQ�<��CF�tц�� ¢�B@Q�<�eG��T��H4X)�`i��i�<I����S@hpzqˆ�5x�s�FN�<���C8V�rD���.p����S�<�rl��w��]�4ʜ M�����U�<1p�P*Kb�1������A$S�<���R�1j=��*^0$�$t(���L�<y�O�w� �d ��L'n�2���s�<�wU�w�bf�Z�A��Y��Jq�<)�i�>G��`A	0W,j���Bn�<Q2����$kV�Ѷ�l���d�<I6%Qm�F�BO�?nY[� Ic�<i׫�8s~��,��=
9ˑ��X�<iA�ÐZ����M_���,���AV�<��!�}3�D��.��k"B ���	L�<a�eJ-M�5��MY�$'�A�c(MT�<YӁ�B�R��0ϒ�x ��;dR�<�R�[�䝀�%1�M���SI�<y'��c!���&�^9a����F�<�� �3&�Z<�G�Lb�Z≚E�<!G��Tת����g“�m�C�<�Պ�4_��L0�^�X��ЪE�<Q��[�A~��I��] ��;���h�<� N�d`f�A'�_�ij�	���d�<��G.#<"%�g����9�w�x�<�BO;A��Atd��a����A�z�<	�bQ�v�����eL~�z�,Bi�<���0a����F��P:Ĳ�a�k�<�t���|�䆓TE�̪���J�<�  �s3��T�dH��c[�1����"O�`"ࡐ�t(��1g��c�^d�&"O$�еg�5gڔ�I��\U�z�Xp"O�l�U�O�:��[�٧S{�*@"OBe`%�tr<��E��e��"Of<1��jI|ܙ�n��p&�F"Ofd;P�7Oqh�P�:H�e"O9W�P�p�K�)L���#"Oh8	���S��(�LBȆ# "O�Xx�fX�} ���
�l�$R�"O�!z�N�+���� �X3y���0U"O ��g	�TF�=����E��9z"O�%&JrT��S˖�7Vr��C"On�b$
�]��lqP�B!6��%�#"O��!@�:� ���ΔSm�}C�"O`tѡ�G	Y��hso\>K��I&"OFs���?b`(HΗQ1�5D�l�A�O����&��>e�6p��$D����Mp�a'�!L2(�*O.�!�F�$(�Y�Eb�\q` K"O�e�0�R4-Y��Z�B?mL�W"OT��C��J��4�ʥa��*c"O�kt@]���t �!E�e⭚7"O��i#	θ(��)�2-��iX
A��"O����쁁��)gL� @�=A6"O
 %�A{8�'+֡}�����"Omb� �'PP}��%�7)&���"O(���Gǥu����D=%�I�"O�ِ��K�2슀I%���"O ���� vޥ��C�6T���"O�q�B���tZ����l%jCeq�"O��y"�ɤ\x��p�@�K��t"O�aꠤ��a&8 b!�)�"�"O�����|�������$LH��7G@<�Űw)
+O�\H�>E���/iH��F%ڑo��D��H�y���:hU��L�)�'@V��B��ќ�ܹ�Rl@~1�pΓ�?���ݛ-�6���O�˧n_6��/�Ũ��w�	�����@�pl�A��}֜��S�s��O9�Xa�@�)9���PZ�F��ѻ��x�Q���<�}�E�4*���zbgH9Ek2aҷ��[y�[�`�<E�ԧ[u*nbr���u��k$o��?Y�O�c��'�� nl�i���ڸA�th۰�ېW��X�q�<١M�>� ÒC>	�O�,�$�:���嬴�v�O� �''��
ӓ-�xVl�1th���=�n-�g�1Ol��%&�)@���"N̪e!��ճ#�B�ӓ"Q:/�!C4���'!�$	�+j���.��+� 	* "��%	!���)���J��'Ƙ�:堔�*�!���}�`���n�\`����"	�k�!�F7=��K$J	
cBT!��U!9rh���S>a�B0�P����Ț{/�"��j��	�'�f�ź��T>Qc_>5���_���"��B��"�
^�L�,��D1D���
_w�$!��S��t�9�'��zE���y���A�'z�����z�՘��^>�CS.D�s�.��&g�@��b�G�4�@ 27�B/;�*mzF*�+'z��)� s��Y���&�BL���M�/8����_�4]�B�<m�x��O{�>U��CU��{ABϩ	��r��E�?�dX� �8%���`)_�<E�DfV�v��|���b�<b&E�7	ed1b�O���'��M��ӯW��� ���>'�Z��Fb��HOL�2a���Ҹ��OS��b�D~��ye�ڋ]�P�i�O��kD�K���=�ǨB�j@,(�|��1ӥ�}�<Q�ɏxh�d�ŗBz��J�z�<�8���`���d�$�B �J�<Q�P0��T��@��A�h��3�RF�<��69�R�H%kSj�avfX~�<�bJ�#�R���cʹ"m���F'�~�<� ̙y��O?IDR�ȧ�i(dX�"O��঩бU��� i7	����"O8�1 J�?�j��Wɞ�{�й�"OP�5�ŤA���BQ�Х$�8)�"O��I����*�W�Ůb��LKc�PM�<����YP�K0j�*X�(��N�H�<��A2O�Ѐ�2e�R�8��X�<ID�ԎO0� � C�&����W�<�)�?���ta��������Z�<Q�g�%5�h�h0�[���q��&QB�<	��O/b�� � ��,)�L�0�{�<�Roȓ ����OD(<�vqT!�p�<�V��s�ZaC�&W:?qȸ{R R�<e�5'��s�	�3"�X�S�dMT�<��d�'*�Aۡj��p�hH[�Xi�<�Tn�
��5��i��xF��%�Hc�<y4�I�^X����E4�({�o_e�<���G�#��j����}��(h�^�<I�GK'{�<p�M�� ����Ň�O�<a"ȓf��k���@��Ta��O�<ٵJ�T�,)�1$��,l��iAI�<�݈w�LJ�H�h�
TG,�i�<I���"n�Yס>~B��$�a�<)�DD;O�@��k
7g��(yAe�`�<�R��K.����+9��e�D�x�<�� ��9
P�ԤB�{��#��u�<�$kX�*J0$�����sh���l�l�<�AI��<.�%���>�d�@eQ�<�я��Y���+w�Γz����ly�<I���#�~�bPB��v9��ot�<��j%W�>	 rb�G��:W� x�<����}���q�@�r��^{�<9��?B�<9�����TL���¨�s�<��U�[�r"�!A�p\����&Dn�<�F)YYC�@��
S-wY����t�<qb� �N@���@�A�
 �ѣBx�<��D�2x��um��No�ai��k�<��J�4K���� -��w�
��Ѫ[�<	���^?`)9T#�"S�H����Y�<Y��فb��t���Mfr�IE�}�<IG� �U��͒���?@��x�P�P{�<��N��%l�۰D?q��x�c͝p�<���GX<��G�f����@Ut�<��jP�����ŅTP,�@�p�<�TΉPC�FR6?a��b��Zf�<��c�r��89��׭
��	Vb�<���UL%p��ݩo��A�f�V�<Y���)$��IG�M$P�x��	V�<�Sm�-a`jŊD\�\JirCM�P�<U&�<(l�@�&)H���  ��M�<��j��֣O�o@@�iT'	^�<	R ��~�� r2W6I�b���̚\�<A�c�,{R�׽^(�I�n�@�<A���RL�8��!V J��C䉁���o0���J4�
zF�C�I67�J�ZsNF�Z�����8�0C��#[{6زGF�@�y��̒�vq�B䉴�^� 7�δaO�abVE�5k�B�I6֊�1��~���u��?��C䉍a���Gx�%��D.,��C�I 
9b�Js�M�Ą��q��*0%�C�ɢj��'��V�V���M�Y(fC�ɡy�8�(@�]�B�,��g�
}�B�{t �a�>"�I�`Ά�v<B�)� �I��NA�D�Lt���(2|�K�"O|$W�^������#M(*�Ũ�"O����j������-�D9HQ"O�c���+Nȱ�L�==��9T"Oh�p���/r׺�c�F�=�͈v"O�m�aE(|�p5eE�XX�i��"O>a�EaP�"�D�l����d"O,$zb"G��Љ�m��JØ��3"OpK�`]�2~���6�5[�,��"O�E/�^/LQ0�'���`�"O��F�ܪ5iT1y�H�V(&Л�"O����3=`
Y�e�f�:��f"O|�t�X�ۮ4ڱ��0��eyq"O���ŉ��k���IՄ�$(��=�E"OXy.��\q��B�	J�bz�4�#"O�����k��j��[pP)�"OH�C�4I|@�6o��X��	�"O8���I��PH8�'����(d"O&�з�F�H,�(�(��q��ٹ�"O2}�񋊔c:T���(�~��5�"O2�*�ߕNʶɵ�O���q�"O�x: �YJ!��0�)]^��Xۄ"ON	!���1M��(j@2\�h�K�"O�}@wN��E��ʔ�L�[�9�"O��Ks�ȗ"��+�J�r��|
�"O\��b�c��27mB&^K2$`�"O�tbT�g�0QǫÚ_H�3"O4�@�N$Dh�� �
W���"O�0�J�Sf��c��^�铷"O^a���EcD��@	R�f*�4"O�;R�G c],8���O��� ��"O��1 'I�}�lm�aAML����"O=80��+Ш�r��R
B
P`�"O���`MM'Q�
�#�n��b,&L �"OH��Q3YyTuS��_6\)�X��"O<mX�)�:,c��{� [X��t��"Ob}+உ�1�~0 @�R���J "O����MT�ǐ�QE�Q���̉�"O�U����-EY^I-ѭt*$H�"OJ�#��8+:}�0n!y&�D�Q"O���#�6m�8���ؿR�0��"Ozݡ��ZzDH �C�k�v��"O���ГC�����B=+T�\��"OZ�*&�Ɇt�d��a�9>M�t"O\���/�92-4�q`��2[D���"O���1��~=@)O_�vT���6"O` c�ְQ���sÆkN(�6"Op��"��V{^����/c
P�"Ol��'�;d�{�ia�*"On��.Wx}P�[s��z�����"O�-��DŘ~��`�T��2�� �@"O���K�1^l��
�{�<�H�"Oڰ�5Ɨ52*��@炖cbx��5"O�U�pD6k��]!��DPa�"O�y��gҥ,�F�O�az#�"O��)�$�"�y�R5[]Z�A&"O���z�z�H��$l|Hh�"O�Y@獟�r�B Cd͙�#O�:"O�t��D��R�)S�+��C��# "O̝@!� A��l���̜!�"ODQp�ъ���Ѭ��I�8I�5"O�ѵ��|�T	��W�l���'*O-�C�,{�=I"��hW
���'{��&��t�"��P�p�J��� �A�d6R_$�b��5g>�x�R"O�=�k<byBF�O> �"Ont r��iφ*�%�t ��Q"O�����#P�\p���i�hC�"O4Y����@ꦇ�_�|��3�Gl�<a�m�5Z\m�v�ʳM
��PA@�<q@LT4M��������=tu4"�~�<g�	U�z�Cҟ(T@TC�{�<Icd��_���@K�C�z]`vd�c�<I�j�V�x���H׼9����È�_�<�%��KO쑢fZ�M:V谑nLT�<y�� ) �xq္�$�
�P�<��Dpz�ذ�X!�gaTO�<�D	a�`]��˭]��(�@�E�<Y[�� �w��/q�I��	�P4
B�I�n�Z��u�P�r�	#�� ��C�I�9�h�c�������3$_�C�	7f)�E�wf�H���{���,�ZC�	�1�P1$@&Z�U�׎B�]�$C䉐?@��aD�	��I1B+��T>C�I�v���H��2]��h6ˊ�6C�I�
�6���8c��!��#���B�.I��4�U�XQJ�(֧�4"r�B�	��}���~f��c�Bb�B�	�)����@ZcF���FZ��B��7���s����=i�a���B	O��C䉃B
�Q�js������C�	���t�p'
�7�����p�C��=S".����I�y�`bW(�^C�I-���p����$�T�vN�B�I�}r�Dra���/�l]��Q":�zB�Ʉ/<x�S啧/��ãN��B䉉2N�r�^?P�~�`狇�:IB䉑/^�B��[�\x��cf�C䉬W�^�c#aU�)�8�3>_��C��0=x ��GÎ5
�i���1ȗ"O�Pr��Ryv��ҕM	�1�DZ�"O�$#f�͇E�+��3g.t٤"OT�#����*�Ȁ�6�L��"O�=z%LϿ{����D�ęP)�"O4mKӡ�/�p09�ė�8�N!��"O�� �+[G������iX�"Oh�� +�F��[�����`�"Op��Eo��^fl|K�^�y�JI�"O�(��;k�����Cm�}��"O��`��S�ʹ���*TW<0�"O�Q�q�A93�@y�"��e��a2�"OƈH��8 掌��%��b�Ry�"O�a�*@�[jT"����}j�"O�� �&�#)�(�H��M�J8�4�f"O&��HĹJ��m�ǆ�!>H3w"O��cn5Z�AhR@��GZ���"O&�y	�LP���I�/	��j�"O��`M�L�P �]6gҾI�"O�	�l�������: �i�"O�Q���r�����  �"A"ON�;LP\� �[F���j�08"O2l��j�`Ԡ��ǘ�@�k�"O��	&�ѻ�)�'�<��"Oh��6LF�Z�2�{�蔶<���"O�\9Gn�A q�C,S��A�"O�Q��c,8'����^�}|�hQ"O�����a
��Zo�1�"ON���   �P   �
  �    !  �)  �3  �9  @  pF  �L  �R  6Y  �_  �e  l  Sr  �x  �~  j�   `� u�	����Zv)C�'ll\�0Kz+
�D��8�1m0u��+c���Gl�O$ a� ˊU�:	+����Tʠj��CHx4��>?B�e	�-�;P���kJ������2�%��ėl��9���o�mX��2	}�	6G�X@A�s���<r��)"� ��Gd6���O�Jt����<�[�e��rb�U��N�IYjp�`�Ɵ<����^5-bcJ٘�M#G���?	��?A��?���18���q�HQ�2�h����?Q�����%u����?���R7�����?qbŪ(�bd�K'-���P�ܿ�?y���?����?���?���غ��b�O�$��c�^�!�hZ�hc��2�
�
Qe"=!#��$�(�l�2}��U��j6O�����A�x}��ɨ��={O�,��#�.J@�A�ۋ �I��O���O��d�O�˓�?�/���-�� ͂*&�`a�˒TF�d�����զa�ڴ�?��i��7͝զ�
ٴi��Z� R��`pID)B���D�l��dK �S�?��.�c*�S�)_�[A|���c`����0{�,�[U�L���qٴ@�6�O��i��=,Ρ���L�`���ņR"I�F;��]78i�f`ؼZ���`�0�ۆM�a��!v�ͣG�7�L�AP۴<�QH!�ȃl�$	�"� �v|�P��8�,(���3�/p�PlZ&Q�jT�H2` ���+
� ����/Y�rAѳ�C��B��:�Θ�u/>=��1ܴA�6�n�d���6t`�Ԡ�Y&��wc4���I�-ݶ=�
s�In��5�4�AS�ۈ�D��đ�I�����D��8x����0I3��ǽ1��%�����'���'���IGk�8�`��O(۴��6(�d��dA����i�OH��&k�����O&�S�OF���� x��p_�8Y�iM�E��XY����7Yx� 2�1Od�SݴB�҄{B�ː��$�lӦ01�,�*`ʒ!R>jzaxrŉ!�?�����/�\�BO�('�X��	X�!p�]�4D{������'����g�ҳLy�T��!����?!u�'��Ao�b�f !�57jdٚ����'������If�9 ��6E�>Y+��CL򐍘��#D��x�D2����6r��Af) D����C�4�>q���@c��֥<D���RK�1g���J�Ar�|��+8D��;����$���x�<�Ы9D�(�d��B`��"���PC�$
¦����0��<���Z����	��h�����su!^�CΌ��-N�B��}2�N}e�zg��h�
��e>c� T�O����z�I�	��q�r���Or�M�v3�	S��)7��c�b�)"��XR��F0�0��O�R�ZPNP�y'��z���%ңH��������<A���֟X��E�L>a�D�=I*���P:<F�5�������?������h�ĊL����ߊadp�2��6`���'���?9�R,��|yb\>�	~��D��Q�ʔ�`��<��!I��򤆔,Q�|rL?-.���*�
I����ğ��y�0W�� f�Z��`�4���y��$��d��j��{-�DD�F�y	V#?s��`k�q����C��#�yRcD�R�(tp���n\^��u�N��<1f�ր�?����?qG%Y:r������Hnr9{%���?���+������?���r��y�L��}N��%?�y�oA�ast�["�ƈ�������6�0<�a�ig�Q�A�G4&M�t@+&O8-X�%;���ꑭ�%'��!Z��$�@���g��-m��<�񨇶X�,cO�g�ڄ`ڟ���ğ��	��%?��<����>���0&sVdqcTߟP��	�MCA��uk�h�v��hƴ��sŏ 7f����h� e�t'=���?�;����� ���IS4h�����X�<�!Ņ*J�l5�1��8���-CX�<�f!N1s��M`r�ɲ���"�|�<Y cH��YHs�ͅD�.���G�z�<aED��R�r	:
@�uri0OAr�<�q�
5���'�RTq��[R-R��Ms��?�� T�;a#W��?q���?���տKa�E��LIH!�Մy#HYy�A yP4��K�#u�&�����Y>����CC'f���F+�.P!0���=��q�E0�yb�ؙ3BdB���yBʤ�rIhb�N��!��U��?�_�h�'�O
ЁK|�IԟT�Ӂ�X�Q ��g�ԭ6_�NP�ȓ=���C���o%t4 �Ŷ(��	�'��7�C��e'���?��'W�`��X�j\د1� m"��KY z����ǟ��I����6�uG�'�R=�꽉�++V8Q��lP� �zd��(!���0!2�c��<\
U��ʉ,'�I@�O�	c��ڳ�@̒e�������!�,Nl�K$�O�t�Y�7�t$���]�0�P]�A"O��BC�C> �ɠ�.�v��Н|r�x�ēO���#�q��'����cV�0A ^�℩��'/"ʃ���'��i�)�⠺��z� 4�-vӘ� ��I�!6��)�v�W��m!Tl3�<�0$CE��xr�A+u��*�M�F�&r�|HfoW'h��8�ɏ4Y��#'��]��O
�ѣ�'�R������+���1� 1�d}pb3�d4�O܁A篞+~���ϒ7&��P��'�"��S�j��mz5IKf���`��I�:r_�dp"�ޟL���ĖO��x�3�'�H���0��Mi�-�!�y˟'2�\�̥���_�̡I�ä�,�����)^�=S��Y�E	"7T$�/�#Q����s\�9e��?W�u*�e(�f�x_w^��^>e���9m��*�Jɱ�|]�T�:?�e�Uڟ���P�O��Fq����ݓ�=��(�!�H?N�� � g�7��,!�J�$�џ�8���ϧr;�E�a��P�F�S�-,���'�r:Ot S��ϴs*��'���'��n�	u4�J��P�N��|r뛦����a4P�7��xZ���_טO#�'���Hf�?$�D��#'��W����l�Vx]2A�i�ة`l��>⺓�D�1c���HC�t��`�e��m�R`!Cr������O���:ړj���`7��!�Ń�������'J��@���r
N�z6�z���+O6�Gz�O��^�0�@K/<���t�РR�b��H㟌e�Aɟ��I�p��/�u��'�B�'�ؤ�����0���vh۰k���ƣ^�t:��Q�f�ժPU4�D~b�^t ͚我�����C��0p�����A�MQa�ܦAI�3��?<�U���ߎ!��'9�U�'.!���"���4(e	ã��?QU�ir"=A�����RY�Wʛ,SI�f��s~R]�${�4�?Y���}�Ԥ�>��w����\i�`I^���v��[y��'6�7��O�ʓf��̀a\?��ɸx� ��Ɖ��V'f XF��92h���ޟ���FƟ��I�|R4ڒo� �iE�ʤ̼�D��= ��R���a���E�7m��Щ���C����1Br�҇B�'�teB��_�=K��@�#���R��&!LA��4KQb�	͟��'{@a)w��8���u~�8{J>��c��b3IV�d�(5K�2@�`������?1'A�z�� A��7:��2G���З'&�0(#�|Ӻ��O
ʧ44k�~	uh�]�t���孉$W4	;���?�AB�h�F��A$!c��A�Q.v��k�deH(W��(�ָ,�����<d��'�B�B��NL��8��Ƶe���%t�M��O^��hW�Z��E��D���[�-?��i��]���`D�$7Ob]�:
Va⥯Y�u��I "O����S�!a�EH�$5z�@Y��I�h��L��%\�7V��fR�AX��lӺ���O��8h�Ph��O����O��di�Q��$)u� �p�'�`R��	-�{�	F�p-T����chb>c�L"���~Qz��5́gX8 %�4&L��T��h�(uC��e�^b>c��i��ёCȦ��	��x�#%Mަ�!*O�q���'��t�OM�OѸ 㖱l�Q�nT�A�����)D��X���D�<�cOTqo���'h�<��	��M���$<�� r�F��4���N��F�ɤ6e,��D�^�C���F�&uQ��&2<!�D�3n%�-<�}�e���M6!���T� 2�j�Rq� �ɺ>4!��&�:t���Li3������'63!�dط���"'+��=.J�`-�#'�}����~r��8�"��T�̩Ta��'I'�yR��3s�� @ƅ�0 P�д���y�DH�du2a��^�дhB �y2��d���j:��)�M���y�&P���Ț�7�����	/�y��\*~�J B���oY�ղ�� �hOz�`�S�(�$�#�.K1Gq���
NA��B�.zB��R�ĮI��$�G�?̂B剺?�$���H�/h����<!�Q�r��! ^�>���)�0F!��.,�5���R�s�P�(&Ƈ0�!�dP�( ����S�Y�����(�r�M$�O?�`s��N">�C��̛0:t��'b�|�<�	�S��}{�`HT��%��c�a�<y��Ȕ\z�%�KZ'QLł��Z�<��N�#,ў��f��9%�xx��+�S�<!��
�Al<�pHut�`�#^V�<�@l�
��Da�ݙî�Z���Uy�[�p>)�#�51���IrFю$�q��N�<� n5i�H'���'�B3�,�3�"ONиe&� u���'$4}�"1:r"O��'Ȭ5n�Ѫ�"_ ��H�5"O8pC���k��Q��R�r��[v�']��'�Ƞ3�lJ�#B�A!-©p��)��'�xM!��9	��@�P�ػa�t���'��Hj�Ǝ��
B��.��D��'��}��掛O��{��.5��D�
�'��Dٱ���PY�E��:\����'�"��DNnx��ۃ�� ��S���F7�Q?�c$�&S'JA�vI���E�5D��I�� =�B	БgQ'E���bA)7D�PS�3,50l0j��~� <�F
#D� �H�T�baT"R�@�.d�"/D��S�N.-7,��T�H��BJ,D�0�T��� �6Q3V��%��A�F��O�����)�'W�yun�k(Xl���:�� �'*��%�rid�
VEPV��
�'�z�{���+Ҭ6�nء�'W �X��ױ$
��2*W�wZd��'n�L��n��>�sb�U��tl��'BV%���5 %���;{���,O�iK��'|�@h˞Pr�!��ƀ~��)�'#�"���M��axfJE�e ��'�
�!�#ܢq��m
6{�th�'���P��,{�Hq��NO\�"�[�'6Vͪ�
�46��)p6�ӓO��m��0B$���R�fɰ�G�!_�t���n����~8�xyG
H�.�!��MU=OA|���
׼�G��)I'n%�O�w1��ȓ-�X���-Ī(~��p�T�]���ȓ �j�"��)�� ��ll��ȓU�������(�Fyh�i�eD4�F{"��ͨ�܈q�8��&�WӞ�A"O��1р��4㔠�&T>ˈ�p�"OR+WHMj��H+�	�!�F���"O�Ir B�%���h�畺:6��E"O�x"'�o� 	���
#40�`
"O�D�$m<#
)0��H F` ;��'-�=ȍ��J�<!Zc�����i��3sjU�ȓk댱�Pf�R�jf+�/�R�ȓ�U�C�Qt�  �-��%t@��ȓ"�v�!�K�,vy|z�	�1X��ȓ@��9��ߡ"z��B��D�Յ�K����i����sR��
@��'��Q�	�-h�Ũs�S��k�c\ Jx�نȓPJ�ځ�8!,N��ChD1;�b���MZ�)�(ʹz
��ad��Z�BI�� �~�4i�A9Vqy7m��R�b�ȓ[���EӞj�x�b5�����I�o?����Q����ƯY8Z�D9�Ǻl�B�	�D�n!2��=i�:}�F�J�1�C�	<NVa��D�C:XU�
�j@�C��8�
�j��@�G�B����,-��B�"%�����A�e�����Y��>B� Y��˰ǆ!���s�d�X� �=�ׯ�F�Ok�M�.�.l`"��Z��l�',�z1+��V'��	 M2i��'8�$�/y�D��@�=�1�'CT�A�F]!j�&�� `߿7>Q��'�4�	!�P���◢)��1��'����Y�J��������MF����u�bHEx����doJ5r��A+_��c�Dұg�
C�	;\S�19�M!s�����ϵP�B�)� b��j��A���y�FL����"O:�c�eM�f�֡�g�ЬL늨�S"Oڈ���⤊�!Ѓ[mf�1�"O`=3��[3st-zAa�~d��Z�P��+B:�O� !@*�L	9�Z�cT�	R�"OT<���S�Z�px���CP!�W"Oj�i��Ǝ3���V����L`"O��@ሃ�=$��P�Lש^ybe�"O8XPGދv����2� ]�"<�a�'t�� �'�v(��B��ؙ��ʫ3hd��'l���QF̆[��(���$}@���'Q� �B���,Z�������'(��c��^8t�>"�����f���'��ȆO^^����"�ͫ�'`��d�*ڂ0p�IF���x`��d�'�Q?	#bAR����G��>8�i%�;D��(���.p�1(�o��²գ#l9D�h��nY!͊�I0E� X�)�q�)D���T��@W�Љ�K*<$��"D�H
��A=a��D΀D���$D��Ç��=4T�!G�r!Q���OЁ+��)�tV`b�ꊲK��Ő��ԁ["���'�B�b�3��i�͕�K5�!��'
�	���V�z�2�h�t/�L�'�<���Z
j�&�0������P�'�ph�Ƥ�&�~�;��ʚ7	JY+�'y$@KAN����"T�
�/	��y*O��	0�'�ڔ��&�$	�:��J4(����	�'@ʀ��Ʀ3��`W'ђ?��Y�'�8r�T�u��u�#�-N���'6�(C��}]�%"À9N��Y�'�HI1�H�/:��=1�ax5�������\R2A��NE�Dy*a����:y"T�ȓ$z�(�%MG19�.@���-Xr2E�ȓ|0���T��s�"�,zLd���M�����CpŶYfC��	��i��F[aq�kK+\�L�x�%����8��uBT� o����3��!0�aG{r�B�ꨟ��A&�&"Ī�B��I�{��c"O�]P��C -�\���Q�̅�$"O��ą�B4ۦ`��]����"O0� �`�!t�<a�nؘP��]�p"O�Hy�S>?��D��n3�p�"O�}x7 �+O0u1�.�;6�9��'�\@���� G!�R��+�����R�LYՅ�R�P-P��8�����?i��х�c���!�N	->e)#H۱z.�ąȓj�t���G?	�*XQ��NF$}��'�P���/^�*���K��a��9zJ����'��5�炿:*4�'a�a�	��Th�V��U����� =s&Մ�I�<8�39���X����vr6�����	#��1>$\u �@E�kRBĆ�U1~q��=}�~-P"��,o�B������F�aRڙ����r����,a���#_��C����P@��j��C�I=�>����H8E��В�%H"��B�I9J�~��"N�O��P��j��p�B䉬��S�ҾJi������	ӊB�ɯXК�a4"߀V�h���+svB�	�k��4�an�<�N)q��63F�=9�U�O��B6D��X�����e�5u�XL��'���0`KH�9�"%��]eB���'A(@�]1�=q�J]R
\���� ����L�!�倚���C�"O.xgѣHzvբReH=D�P���"O.͡��#$�QÃ�D%\Y���b�'���ɏ��S
l��|���\
y�.ڷ1�H݄�0�(�qf��\p�����J��ȓ~hz9 %�M0�uK�ܕTm�@��@�\�s7�
�L20�!E򢉅ȓl�y�Gm��.Xɂ��Eo�\��.z��œ�Dʗ�h�pH�'����
����RWo6I3GkZ�?��ȓS�$h���Z�|p���L	\��(�ȓG�\�p�H�2�\؅�.7�bl�ȓ<�졘ĮҰt���[��(T� ���W���KC���H��#¢H$L���	7۲�	�Y^�9�4U#�-w#�K�C䉢H�va�%ŔBz���(9��C�ɆQWʌ;V�_%=4*R$OC94Q�C�ɋ^q�5a떙C��@���VjC䉴tֱ�جY~��Ս�s%0���x��`����^��������Z�F{���ި���A��&�P"���x�F"O�hR&��<P����"O�̒�!m)\D��e����2�"O�DyЧ�3@��\ ��%�L�Y`"OFXkƠQ6l!������x��Ĩt"OD5�s�J�b�d��G�Ȩ;�`���'�R�Љ��Ӊl|���`�4ƀXs��Dx&Ն�k��{#�Y���L���)լ��ȓ �$�󓩍�mT�ũ��
.�le�ȓb��Y���CX"�s�F���J��ʓV��rVe�61�Й�o]0i�VC�I'�8$���A3e�0���7Wnbu�=P�k}⃚7Ŗ��J�O�<}�b� �[�����-�� m>���\c�=0��?	��5�⭊ƀ�d�ܝ�$���mZ�O�y�o�3.��ˌQY�퀊�D;ui �x7C��!ɮ)�#��ć��X�Q�JT1f����͗ˈO����?ъ�� V�<D�D	�t+��ٔ����$3�O���E�+/[���@X�>����'}��5m�	��#�"g�t�t ����`�' �ӳ�'cB�'`�S:B����	Ɵ�����L����i�9s�D	���UԟI/y�f �N�	*6���ܴ���y�'
�@RD�WT�^ЩN܈��m���9����T�#͊�M����")9`����CU�:X�w�V9KU�0e���y˃%�?�����4���@�K� \r�s$%�
�T�L$D��J��ݟV��qX�A�'�8F=ў[��ɝ!��E�Mޜ'����ꋚ5���O���̋C�Zݡ$@�O��D�O��$럶���|"`C���?�rdp3(�[1.I R��劣P); FY!`)�|���䏶p�,�@�m�[���D�,O�<�B�-~�\�	K�Xǐădm:�D���D�,Of9т8s�՘�/���nPqҘ�T�1��O���7ړ�yr!�r��9Ag+kH�����y�#�L��H`�ŝ!-�|ٗ"��?9��i>5��Py�.��	� |����6Q���!��y���!�
��'^�'F���'�3��% ��M�e��2o�+4�0p���%�~��rE���N	CR)ϛ'�8G~�N�
@�H�,�..���A�3�>��uL��"H�fO8-�P9�)n�D7-�k��R���\��Y+D�D"f�$A����,ړ��OpLJa
 7x��x"0Bh�LU "O�t˖%�7@��X����~9��gR��ٴ�?9)OnM�!�H�T�'��M0s)�$�5�J�:Z�i�d*�.2�m�\���'�r��+I�(`��F�?(ٚ�D���;_[�m�u�V�@���J�	�,@M�TE|⎆/YҲY2p�րo��A�nĀ*�j֝�B)8���ի1�f���2�f�l��' ��Ο��|�U�j�*$���X��qK�Ey��'4QS��d�8ȡ�ϡ9���k�Fw�I<�Z,�qZ�1���A��5�j�Y��?y����)�|�L�d�O��S�̀�J��jAM�"&�`�&�O,��',��!��)��gL�"��B�����IV�f'ڽI�eG�EFp�"�D��^6�|Z���nT�Ie�V'�;�u��.�I�;XL	��BAJ�z�̕W!�$Tp?���������� �0�f[�p���h׈��t�2)#"O|�3�d͑qLr`�4��1{T(���I��ȟ� ���E�A�L)�z��v��OZ�d�O����
�$�O���Ov���O�5�ThH�e��IчB�>p�ތ��C|�(5(]�}\FUr@n;��'��O�E��Kט	]�-�A�M7q>.5P�cS��5��e��"���֣P&I�)�Mش(��ɘZJ �8a��6����"&�3sgp�n���OR�=q�'V`�2�W;:�d����L���!	�'/� Y`
X�%N��P)�������zY���ҟ�'ij�zр#u��0���
8h �x�bַ*���I��'�"�'�O�B�'�	�&�Sv��'0�)@hE���@ġ�EJ�A��N�̜�r�W�'�Z�Q�7X܈e��Q�N)�`�ۀ;��%�!�AbJ�P̘�8�v7M^/VN����Ū�O�� � 0?NJ��g�M�p���q���O �=���DÄ>�@��#T1|�@�q���o*!�$��xWlq�ڵئ$�1%�ɇ�M����D�9XN맳?ٙ'�PX��%Ҧ>z����n� ��:Y�eb���?I�(Ў��`cV.H�R�#J�	�6����p�`"{Q������LC�! �$Z��0g��'����E�M�`��M�� ��)DM<%���1�J=p׎Ƭ��'��ј���?ٍ����'>G�� ʃ�twH����"��D �O���6㜐���Q�$XD��岷�':�%q�T�� z�v��b���2�"�'R�'�B�i�O�才<pt]cs$��.X��W,2���	�#��%#�{b�	
d^��n�:*D"�9VD�[l�㟼n�d��	"��O�}�0�@����հoWp�#�f~��DޗyC8�IyD*�$�O����O��ɽN�xq�A�}V̸e�!S�����Ҧ����lU���<��H|nzݕ8Οklָ5{� �a�P�|ISEj��0<n�����?UHנ�y"��H���O,�)�O��	��LA�ģm��%82��0&T,lСn�O��DX!���b�Dq!l�?7��)5���U�G'|�,�HOa����Y�x���ߟ��
���I�Ob��蟈����}��84�V�0Q,m�R���%���GR��$�O0�`"�O�	(4P��s��Nĺ����R8�"�U�����hKŦ%�b�R��ߟd� �<���?a�'���%�Y.�"�OE5���k0����yB����?i�3�n�OF��>��s�b�Qg!H0?h0�q4d>=,�c��s�oZ�<��Ç��MK�iA��y�1O��]�?���aɀqC/A�1�֑�V ��}��4o���c�'�Da��?Y�'�?)�'%�O�8k%m@$�~8�V�B��M���{�0]c`��O�˓�?i�S�g}��F�b~ 8e [U[.1z%F�*�yr�ݑ2�9Ć��FϨ�3��Ͽ�M[����^c�SLy�]>1)��ͧw��}١�F�s����H����)�"�S��.ڨF7�+r&�#lD(������'*�'�Q��K憕�a�Ȩ7$kh�c�&0D�d�P,Q/BtD$"�n��B)�\$,0D��k�M��AE48C��TY��%;D�X�w��ZvE��!+Y�p�QM-D�(;��B+A|�b�㜙=;�h���&D��[�I�`����s_�V�!��$D��{�	�1	�e���P�'J����=D��`�Äc܌	#1n�+ԸPq�(D�ȋ5��=�(��ʖQ��Drp''D����H2b'n�E!G�-<ā�	(D�h�6�*a0t���V��s� &D�P��N�`/h������`�$���u0^�!�B�E>��ȑ��	(��GbW>���/ZV!�y����?m�y˧m�����UC��v��s�̒�J��I*QbI|����!Q���
$j�?�*%��!�WN��3'%p�AqDA��+6�)Х�Y?o�����Ov�2Aĕ�g,8P��D�z��'C.5F|7��K[���ӭ�*!q��Y �X�*���ß���P2��=�ԭ��{7`��شd'�X�t
�
8���c�!{�N����4��k��9����Z��5Z�aR�MC1�޼�Zi�ڟ䬀/��p0*af�%Q���H�xB��!�?Q���h�P6M1�L�*q'&ɪ���
�P.!�ոMN�ɲ�G��\&P�u�Ǔ&	Q�{Q!L�e����3��>*t.�����0�?Q���䓗�O��s̏c�}�A	��x����v"O�9���7�X=���� <oa�"OЬ2��]Q8���F��]�I"O 5#��B�lBG�ޥ�¬�"Or(��aS�S��=J�@��4��e"O,��%oǌ H�0i$�����"O����,]��|�
�f6�i��"O� ���
�K��1 �3/0�:�"O�������ы�
Y+���"O�%+dꇓIx��G�Bk:�25"O���)�$�Ls��Ʊ)^�QB�"On�	ӄ��8�g=���"O*�B*��S���g��q<�� "O��K'�K'��-2�XI�U�D"O��a�iҥ_�2D�&�8sp"O�i!�V<)p����dS�I�.P��"Of���)��#
a��BP3d���@"OB8�ՏY���C6��ApJ\I"O�}�Mή8m���q���Y_��"O4��a\�?��5��F3vI.,�7"OԔ g���u����iE�ʑ"O*�(0�Y=q��p��M�J0:��"O�x�s�/g�,¤�J����"Ob� �.�:iB�d��	[�']�s"OLlaF����*?��IIWm��!�D�c�4)6�&*���3բђ*�!�dW&v��m��N/�ʶ���!��9VF�<����A%f�8¯TS�!�4aF m2��4����@s�!�$բN��$
�.h��E2L�!�D
�GJ�k�Wp�5iB�B�!��N�=��-��)�Be� �g�Y�!�dZ�^t�k��|�q'��6!��D?"MDMs�jŕ����l ZY!�$�iV���&�� urb\i��[;/r!�\�M�|$�d��V�KQ��(�!�d�W� 4A��J�H��(3Ӆ�*H�!�䀿O1P)���܌ds�0����V4!��xi�( � Ti�I"iFx!�$�).�P�aë\�HN�������!��
�~ԨUm�	������O(!�$ dC�D	%E��oZ����	Q!��"Τ����ƻ6����0�!��22E� ��Kݢs]la��2�!��_�y^���B��"v=j�Xl��s�!���a�;DHHI;8c+�?�!��� SJ�4懐e4�e��#�8�!��?�ܴ�W��2?�1×Bkp!��? P<Ȧ	��w��1��AL7kR!�T+X��̣���dtā
uC��|�!�D^�~��0:�j�!Y�Ӕ#�* h!�D�(r*�8H�*��G,���
�2e!�DN�hBFl�`	Calp1��	?:�!�D��rB �4��G����L):�!�ȑ[Ǣ ���V()��кV�7�!�D�7�LbW��n��DuC�U�!��>�B���K1]^���b՚	�!�ޞr�~8�aʵ�  �a(q�!�dUF�,��� �4	�A(k�!��V�4:��DG׊=��`<5!�><H�Ĺaʬl;3`�v)!�$ =�A@TFK�y�J�!@ШUv!�.�^H	�KЊ[�2���kP!��@�)>�:�C����L!�$�+.^`��GG��zO��T�!��eN^���HBn�@��ʣ@(!���,R�5��C�VP�6�S�6!�$ܷzN��C�CZ,y��G�&v!�$/Z"�r��<�
�p��p�!򤁚[v�֨'#Dx�2Bj��J�!�D�0�Sv�	)<�^pj�A�!�� �0{ C�X��t��7]>�h�"O�T �fU� �\�pr��&K8�y��"O\�aM�'�$��������U"O����8?��! ��"wf$)�"O,,p�爻-q��Q�}t�BR"O��`V��zd�-�:rxd�A"O�����Zy���`-: �DX7"O�qB��8��,S�+ߌ}�J�t"O�i6�C�KB�J0��	��8��"O ���jJ`�Y+�D��H�"O���#d\�<]L��&�T��"O$e���Tڊ�c�KǟA�M��"OI�f�/Cz�T��Ā�g�D�ps"O�$���.,_� Wc��?,<���"O
�JG��i���`�L��4��|��"O�����0 �M�l�T��"O��K$�ǵ^SL,�e��aY<�"O(%�� �2% Ä<\*�\�A"Ox�R�/��<z��Y�%��l2H�8w"O��rr��0I>�䪓&�2O����"O�A��#�����0��r
�Z"O�ْ�c��2{TP�%�3��%�"Ob��g�B�b����BI��"OT(�2s��rۊj��mw"O�a��ʟ>�t�#�GΐMc"O��s��]��(�&mI/s�����"O��rd"]�HD2��"�T*4�.p8@"O����c���j����N�PxK"O��1���Tq�ڸd�.�ۀb=D��Y�J%?� A� M�B$�X��@'D��6��,��B��s��id!)D�X*aNZ�AF�MBA�] �8��a;D�8�@�=*0�Q����Y@�	��3D����*T���ᷣ�:�ȁ�<D���  �hvvوs��M ����;D�tb�P��X��BO��d��*Q�9D�(ч�ԡ,M�%�4�Ӛ�[�*6D���TgƊy�8��HQ-<;ީ8v&5D��䈊���=�g��K�h��o.D�4�'%Z�mY
���=>Q�1�.D���H���M#�hK�Xb:�a�#,D�Y��7[btAS�I�1��wM)D���1	�������f2���(D��*Be�Lm�rRj�p ��&D��p�M;w,��d�[<6�fe%D����G`����Q�"p��8D�0�\�D�D���T�V��ȣ�f6D�
ŀ�$�ġ�Q*$A��8Y`�6D�<��k��Ml�����Y'
u�L�R�(D����!��\0��ba�ױ q�����9D����jP@�]� ��z��ib��7D�@!biʒG�^���S�O�Y8Ҥ'D�l��C��z�B��R�Hx�3�,'D��YB�֒@�x�)�<40"P�$D��iaR,I�d�RԢ��s7j�h�-D��0B�ŜT�0x�"E94:-��%D��2�a	s�b�XaA�k�6u�K%D�S��T�9j2�q'��0�ꤻ� #D�����a�l���R+k^���1*=D����;���K�	��� �:D��V���%څ��2sO�4˖K9D�P�w�Y�cilQ�(Z�S/fL�TC2D�xDlȎ~XHB��Խ48��;D���U��E*��R�B$
�	W�8D�� (��D�<�N�Q�.5�钇"O@���T�Wqشz2���vye"O�݀�o]FB^�(��B�FF��ȁ"O�!���57��k@A�c8���"O8���`��k��Y��I `Nu£"O~�q��q!����!��w6��"OX1�B�� h��H����(b,��"O�`*�B�I,5�'e�1&��p"O �i�,�9�x]*�V!$���t"O�]���҇�%��&��iJ"Op�+̳hŲ]����=m�Ԁ�r"OΌ1c�,qHE@`�/�E��"O2�A�l�d�n]c��6�|ٓ�"OY�1��:RTf�3v�^p���"O�Œ�&�v�b��ق7��a�"O��Z���G�nqꠁÊA@�"OP3��΢o�H�Psf�Mm<�aE"O���T�Y6<_
�f���aL�!��V��f��Q��n�@���NX�!�_a3t%�Η���9�a�,�!�M�A��X�2���u@����!��N {1h!f���K=����aԭU�!�򸘳�?&�����t��u��8@����	MV�zMKB�˘uc^��(V���A0a��mqo�:>&x��d[,8Y���|������9Q�R,��gP,�
ӂ ��@3��,iVE�ȓu�`8�1&�lY�c2�)"���ȓ:�FdXB
Q�~��F� z���|l��6'��Uh���W.NC�	I����셑9ti#���Vb|B�\�=0�LIW4U�*�+[�C�I�b{X���c�I����6�C�	�Yޔij1*�?W�}�`��w�:B䉳XS�Ah�O�
_U�}�F�<� B�I���y�@��S>��
���r��C�	�kp$�S��zt!RI�C��C�	�E�Pt�e�] Q�`����ǋ=��C�ɥs�غ�i�'M^�W�H�6C�I(q��`R�%��DmaajD4LP8C�	�O��ҵ��'!�:�hV�]�y_�C䉆p��DCі��4���Y�V��C�	Z����т6xހ��mX�p�rC�� IX��SD�ƂYo��C�e�$R�C��)�N �������(s��om�B��;c�>�)Ffc�`CB��W�B�ɑ@��NW�,�3.ɤs��C�ɒ0���� �5N:�X!��H/$96C�0)�׆�B���{�
�1/�C�I�}d���^
hd�2*�(pðC�x�(Qrf�[�e^jI�ƒ�d�TC�9)�lIcG�-�@�8PcF,G�HC��z$h4� /�5c�Q���E4�B�	3� 1�͆?Y�x'dE	��C�	gZ�8�ͣ���v�X�p�C��6*N^ @�c��(���Ѻ7{"B�I1@����fAz��Y��N)e*�B䉽�l�:�L 괔�&�C�ɦ~1��
7_v��ÂW�4pC��J�L`S!̜�|Zh�3�7�XC�	�'�iSBC�6 ���z��W�pwNC�	�jJ`��P�y�����J�8,C䉣@	��c��Cq��9�G�H��9��?V�	;�S�C=d-��	%��1H�v
A7�Ҳ`NB�)� V\BF��Vx�i�E� ^&h�2"O`ܘ��*��g�63���"O|�3�^x�ÅH�![���RV"O ��G��"��fO:`���"O.�X�e L��u��ڞ2�HD(q"O^]�e���g��_�����"O�؀�	��=R`q�S�/G�0�ٵ"O�$r��_�]��	���&�<EV"Od�TB�#H��5E�"]�  k�"Oz����[9=�D�8�䚈��1�d"O�͒O�"F�ة���A�|T�"O�Sa�+<؜�فQ�/
Z< "OR)3��[�/�tK"��Eהd�E"O,��$K�iQ
��&�O�Iպa�%"O ܁���
J��!o�x�.�JV"O�� �Lڭs8B4�(���y�S"O5x���%Dũ��+x�����"O��+�ɔ�S�S���T�"O����#9DΑ{��U�<�>�2"O��7�J#QŰ�կɻ7h,�HF"Oz���/&���K(�����"O�$z�I�,1�le:�L��p=�Je"O$��'Ǯ:��%
��Ѻ4&�QB�"Op���WP�\[EC�'YlL�T"O�����5a�����X>Da�`
w"O`��u�Ӂ}���գ«*2\ "OH`�H�cR������N��L�"O����&�T]�A��e�>q"OAcA��l�(�S�GF��h��"O88��fߣ*b9�ӡ�:�t�;C"O<-��m `���Y�-�fq v"O���ك#Y
�*�A;2�$Uhf"O�#Vxk�tP�BJvp����"O<�G@�6.��@@8o�ɱ�"O4\���c���fj)��"O�����n�x�R�1��j�"O�l)�� l.XcAY�W�IZ%"OL�ۄ�U�]||r"J�!���f"O�I a#9����wJ3	�lAr"O�Z�`I 㒹qר�>zyi��"O ��"�@G����X�}
(|8�"O2%@�ꋲ	P|��f�|�<�[�"O�I�M=:�2�6�I�����"O�@��MX�PڄJ�
ld"Ot�F�I)h~FZ�
Z4�0��S"Ox��/Ӽ:u�!١hď� qi�"O�P�&
I�<Sj8��NS�?B|c�"O8�W��#�`]�`�YOܶɹ�"O�Y���(w���;�L���@���"OH�@�垚$aީ����0�r�i�"O�4x�L#V�Y���#�д"O��b�)��>�h�"�a�\8�"Oj��4&��5�<5�O,Vڶ`9E"O�ԸW��{�aAQ8���:�"Oi�v��/���G�X�S4��F"O�����O6RrE�eB�'08�P"OD��@�*^�M���܋?sZpKA"O���P��Ļ��{Y4 �"O��S�T�q��d�>B� Z�"O��0�͜o�.���
�W�h=��"O�̲gf���s��.� �K�"O���6)յ2�0����G"JP6"O���ͅ�\����
���"O����ϕ�o����xٗ"O� H9�
G�s��CSlͺ2���Р"Oĉ����3��*���x��	A�"O,���P!j���!�:�>�0f"O�(�� ʒ]ӰA3G�ߎ-(Mcw"O0�a��#-�ܥ��g�*M�zC�"O�I�@jB�@�p��GU^� H;W"O�AZTK��71̘�FPn�s�"O�$�,��cVF�nt�*OLQ�V�ʈ^�8�S�,+¤i
�'{��:� �e5�)�hZy���'F��is��T�)�oIY��,�'��0`�EG�0�.��U=9.�*�''|I�p �6rʂ�pAC�9�`�ʓLmp��O�/!�x�p�B?x�H�ȓ
/rI����B]�=���*����v�(���%�D}�4OV�'	C�I&	�8�Ƥ�� ��EI5"f�h�ȓX���B�k@��rU3��Y˾1�ȓBZ`̢@,�Nז�:C�͜E,Ʉ�Al���,�0��T�p>+��l��a�����S� [�Ł�)D�D�ȓ>�"� �\��4�1�U�� �ȓ1���g#��(�
b�Ӝh���ȓ3wP0ᎉ�9��	Õ_�
4�ȓk#|�X�m�*�,Q�BAW/D�V����tiqD��.,���W��v4!��"#D�1�c�Ϟ��C�KͶ?J!���t��B�4?��	�g��)�!򤖳+k��g� ���{@e��(�!�Ӕ5��`�NЧ%��t�e�_ y�!�(d�a�D-���A�n!�ă�P�X}RT�,��ȃ�%�2!��'q�Y� ��UX"A�l(!�߯0�8Y�6���oW��x��S�!�"	��Lq%Ȋ�
Sp}���І/�!���y�A3�ǀ)m����4��0�!��?ɠT��%��60~��`˛�#!��A1ڗC��)�	ѱ�	z!�Č�!@�8�3-�(0�ΐaE	�t�!�$���!Z�*��� �Q�oR)9 !�N=��v(ѺS���:��#!���*�	P)U[CJJ'B̄ȓS��TQ%�
Bi0g��9�>��ȓk&�	� '�Wؔp嬕&\2��ȓȌ ��J<���?�vх�@5 ��P�t�R��C;e-��ȓ��URt`��y�&�1�kۂ}��`�ȓ��x��M����#7eҜ]�JT��w5�J��&p��X0H�A���ȓY	�	f+�o�� ���Cr�ȓ\��6͜;#V@������@�����GHJKwo��\��Y�c�x�ȓ �,Ͱ�Eƛi� 0��17����2���:���ap��QJU�-�t��ȓ=M�E�%�F6'b�Pc�Q�f[΅�ȓ�E�2�?ڐ�'�B	sF
��i ����z�x P�O�D<�i�ȓ��]ɔ�}����+�k����2tS��\2S�X-Ҷ͙8r���R&T��g!ݮ+��8�͐ �8���R:��ͿǨ�xv�U4#������l0T/\'o��l�5�j����pV�ؖ�]-��I!��`/6��ȓ6����Va��)���Bfa�<� ��@!�
�����D)%�iQ`"O��
L@��m�U"��fmM �"O<僲X�J,8A��K�,T��c"O�P���,+ҀKG�0M���"O0�[WF�;\�t0�+E�@��"OP$)�\L�]`Ǆ׽][�}�f"O�麦͎5K���*B
/�b� �"Op�d�,H���b��� �h��"O: ��B�2� L1d"��_��-k�"Ol��Q��I�����>+䘇"O�8r��uU�¡Q%~��""O����+�b��b���|H��"O��z��g����J��R��|�v"O���pV=
fհ�i�!Q�HJ"ON�!��c�D���Hj]�y�"O�d��K�eBDE�`�/^�&��1"O���&N��fsJI�WdEK�$$�$"O@�ņ\O���7Dl�&a�"Oұ���gՂM��
�)���;B"O^��P�N�1��*�Z���"O���d�L$:�l��B/�%lP0""O �
2�۪+F�(A��FxC�i��"OB��ûg�V-q�*��~A����"O��1E!C�W����ࢅ�]�� s"Ob��K�~�r��#$H�*��w"O<[�B��H����e�c�$�e"O�q`�BO�0� rь^��ӧ"O�1��JB�;b��x��% ��q�"O���g�YS���9�|�c�"O�Z��9�D��E��i՘�a�"O�Sg���F������>� �s"OĈ��(�&���T��� �G"O�Ҧe�-ł�в�ɘ>`��$"O.0r���.R �#�J��fo��
�"O��B�E<���Pj�Vd�p�W"O�P7���f�f��$JԤ\��Aq�"O^D���K�w�j�s�ϊ�.K:�2�"O
���ɂBw�}!�ޮ*TH�F"Oa�ᅝ%^��֮¸a�l�3"OƁf���m��c=2��L��"Oı�ċ� ���i����"O8=�ڹT�v�Xu���3�Jqض"O�����"f<x�o��/� �x�"OD�f@кp�z9��H�ZVp"'"Ov�!��U�'�H���*x_�+""O�u�/�`�M�e�I 0R��"O���������R�ˈ�0��(�"O(H�1f�=Sd^5���ʇ+Oj�!�"O�eX"��/B֘�v
�D%���"O2:�#N:�0��aO�!t45[3"O<d�� Q>4�Fa��*�6�%"O�u���L�a�ce'ܷ��E��"OD��F�F�H�h5�1,�#N^Q��"Oj1��K&5}�Y�ԢN1_�x|�q"O��X6B8UƁ������ʥ"O����h&@f��!iF�?��0�"OLe�ǨE+L�Y"�*��X�ȝȰ"Oօ�PK������H�̰�K�"Ob��� �7H-���)u��iR"O�Ҧ
�R�r}�I�T/z|�"O�}�6')yRxar!۶(!�'"O�� �ڈ���3��D��I9�"O�a��i>_+�d�	5&dd�"Oę�t�B�#
ɉ�� �Af"O� ������J�̩�G���e�PQ+d"O����/i��X��ܤB���"O~}�b��G�u��I,��������,�{�jP
�$��%<OZ���\x��m�#�G
"t �b�"ONic��R����O�>[&��6"O
Р@D�d�f�g3z�u��"O��K͐��i� ��(e��S"OƱI��/c���ӥZT�$�2"OR!��&M9C1��'��Q�b"O�l�	��W�1�@���DH�"O�[t�A�>�4����G�B�
���"O��bkL48k~��AT�g뀠�"O�1P�	Q����v�s�l�3R"O�l�2�*9p��q� b�"<�"O�p۷LZ�8�N��%e��o��pE"O�Y�O/W����/V�I��"OD���#2߬uѴ��`O�yp"O�Bcl��7�����09C���W"O��+�LH�m��A�PeH'9�Y��"O����I��`���*K�+z*�e��"O�X�s���#ݔɉ�J�s#�+�"O�Y�c�A^E���hݚx(����"ON�Eɐ&	��<AJ_;7�QBR"O�l)TR6R�"��0��&)���Xc"O��LS-^���Ƈ�xu~�3"O���!��,o�*�A��q�$P�"O��P�N�q#j���B9J:�p5"O�(�&#R�8�����i��`t"O�@J�8sD��;D��\�x��"O8�Ǌ��BJ6�� cR�Y�-�"Om�æړa�"|��ᒇ=�)
w"O�4`�J��XΔ����  � [$"O�`�W��X
L� u�(��"OB�"�d��V�l s���;��m��"O4�	V˗2 ��o�2z���"O\A0F1s%����XUڔ�"O��2�Ǉd�b�R����])ԩ˴"O���b�9�!�aٖV �!�r"O���RˉH.b��Va�43 �kR"O&T�L�I�Bp Baƍ<4�&"O0l��N�ON�Ѱ3!��-p�}�5"O��ql�J=h�Y���.q�Ɉs"O꽠���Hl*b,�#_Bl��"O��cX�C�xQ���,2��Ԉ�'O}ش�A;�ʱ��Kݩ%����'1ܡ���	�� Y�T!��HR�'��9`Q!":���Ub����'㪝s��Ե"x
����B�M�'�$�HSd�5{T%��BO�9�,A�'y
4��-�	�0�R�W0+�0	�'\& 
u'�U���a%  z9�'mޭ���u�$](�C�	�n�y�'�И�U��w�*�{v-�9Y���ȓg�ذ����0� Y�N�,T��S����l{T"Ҷ,�L�ȓ3՚�K�狤���E�l$ՄȓI� ��3 �4�$Y�#%Ibe�Ԅ��P��𤎹�rd���4��ȄȓJ�~}�����&�B8AD"Y#7u�H��u;�m�W�Ӵv�$MHv��ro
-�ȓk\��;�&��H����5�0����ɱņ9(��x�ɗ�^o�p�ȓ�L!{]%��HR���pP^x1V"O����-U�� ��aM�&��6"O� �鹦�ϦN�dى����^d4�E"O���7
ݨVK^a��Յ���x�'D��)�"~!���'�G0��՘�'�������;��KP��>.�U��''.#Q�N�(�<P���
0J���'����Qg�b�ʃ:��p��'���"��:B�`�b�&5��I��'�Ī�OQ8).uiR��4�*ء�'���rHD.����g^(i� (�'k��aeN�54Z�Cp�5 d�K�'[9	7a_�:���7E� �2��ʓMR�Ӄ��/�0� kp����&T�AקÞ9�ݒS�@�� �ȓ/ߢ��! f� dJ�%K�~(�e��"���ۀ&�)d5� 2�cJ�`�, ��]DIJ!Dߪu�&5ÑÉt:�X��X"��$V�)p��"�J�^��܄�6�R��Ĉ �)� 	7�vd�ȓ��d�ɖ�Q󺡰�^���]�ȓnI(�;W�~�<|��5��m�ȓFL�� �R$u����5]���b�����EsP�\����*B��ȓ1��bG���Y��x6�K+;��ȓ(��e���R�8��`�B��=�t؄�-°I��O��Y�eM�S����"���aSo$�r�f�$&�Ĕ����Ae`5-�X�.��
���r��\(%��8X���ѺPȖ%��|��Ӄ��i���b4��z�p�ȓ��c�h]� �`}bg�J�m�PĆȓ�jE�u�C�u5N(:�j�*�M�� ��Q�bO�<^jha�V��2�p)�ȓ`�ؐ	�CP	4h+��ɗ(fD���"Jl�1PdÓ�ܽRG,��ZD��*�:�;��32����5���t�@�ȓ'؎-I�-X-`�"���Q�#@��ȓHx�Q7
���3sf�1:ԁ���`�A�f�l픈Y��6v����ȓY��e3�*O�Mk�����6t�����kw:�X��ͧoi�u;�C̹_z͇�9p���C�Tk=���ĲKԜ�����q�H�</H��B��	B�5��������=��2dJ>uV��ȓ:bft�q
\��ق59-߸̆ȓO><�{Q��i%Ry&�ߟB��ȓH�,pb� � Z�b�?����Y(8���x�,Tv�[*CH��ȓC7����ḳp��a�G��6�^|��1�(�`�� d������
複ʓ:�Ȳ�Ճ6i��� .� ߞC�ɛ`?��j�$5��S���)��C�	%s�Y��Փ*7�@+ +�R1fB�ID�|�:�h�� ^DI4(֫ �*B�	�T��eDէQ�0 i���B�	0e� �D�۠'��zs���B��5s�B4�4nť-��r���^M^C�	��B��#�
D�*�vNݙ\*C�I�0!�ӕc�5@SI�2�[<!gC��=O��؇g�9��ii�#��PZNC�	2bR��tE�,�Z��`�	B�LC��x��wɟ�c�$fם ��B�	�pAr��n�ix%U�*N�C�ɄS�f�;1�[�k4���f��C�ɾZR�S%�����w��=N]pC�)� (���ϷU�HC��
}�Xx��"Odp���p��E)�$�M?`%�!"Op�BFC�+��., d�b"O�}Rd��9E�0d�R�*%~��"O��� ��F��B��4�!�$���p ���{[��"����a+!�X��(�Y�ɱ6T$��׀I��	d��(�����P�
���*��6
P�p�"O���wO)���A��X�W�QA�"OlX	4"�5 �~�Zw �a>�	qw"O����ok2Ti8�O(t��`"O2�C�O< a�Y��ӡM���"O�\��@��<�"J͖x���"O�h��#��(�`G���4�X�p�"O�=���:$�*��NKD�`��D"O69��$�|��U�X��Vȑ�"O��S ��� H�v�
���l0"Ov�+b�D���w��W����3"O��f�' ^��P%�b��s�"O����ΖW�.��TN�/�!�$��e1d)B0��)9�,L C)��!��+CX�x�����A�зk�!�)c~�����q�z(�$�2>!�$�`O,`*!ѷ.tʽ�7Gߐ6�!���'��]+��Xrb%0�&ܦ@�!�D�<v�R���W��&�q�!�D��~�Xp{$�D��4Y�$�R	2�!�Ӡ:,إj��1II�9��KB;!��(h��RU���Tmc�*�;�!�$LQ����!ϳ}��I@��,P!!��G�5^�)�ȓ=+�4�X��P�!�S�Q�����F�#%k�݊��c�!�d��T-Q�I۱ Z,9�b;{�!�J*Qs��`�1p�%Q`6-��򄃯u��P�ⅽ+�8�s7�ʄ�y���~�x��a���v� ��&j©�y"�O�L�:�Q��u�������y��
s��́Wjϴq�:%�����y��Idă0�ܽu��;�A��y�4{�*�!�V�w�T��հ�y�A�A�"	"Of�qR�� -����<Q{���H�a�G�!ȕ��$��xS�-�-i�!+�LȚ$�5�ȓz�t qD�!Kﰨ1��_xH���.H`��þ)�T�R�Z	�x��o!n]��dDL1\Ҁ��)q��� �@zU!D�0!~2��?z-����v���o�*D�,y�w��> �E�ȓ#�h�qEK�nE��⦯�A��=�ȓe,>0{q#0q��Ұ�ϫd2A��a�@�R��G1��]:�L�2wJ0M�ȓ/�����S`y��o��
8��ȓ`	v��� )>~ܹ� ��t��8�ȓ�(Ȁ!G�L-����a��)�ȓEAD���WyjH�ׇ^)A�*���a�t�Ƞ��7/|@j�G Z8�X�ȓX0
�KH(kV�1��}5r1��[��p�CK��
.T��ND��I��
6%�p��N����wF}ֆD��n5j�Si�J�j�b�^C�T�ȓ3��ɥ�� Ӿ�"�A�	�P��1����々�P+��
g&�#�ą��d��y!-K3P��ٵN�tBJ���t@d@kږ8���6�Y��S�? &H�BZ϶��ůˏ f2=b�"OДQs��Z�nc�m�ah<�2"O�xA�X>Ɉ8�w�I<HK2M�"O��q�K�(C�PA��ӝK6���3"OF�y��?1͸	ڳ`Σ���C�"O� y KȡF
R�:�B�n��Y�"OR�i���P�L�cBć 6m�ԘP"O�Ő���< �v�[q�F�G��R"O���D{��AcT�
��:"O��҂��
^����ѽ^)PH1@"OL���kՙJu�� �w���#"O挩rƟ35&��%g׽c�%1�"O�p��(�>1��KԺr����p"OR��7�@�nL#1�5;bht2�"O"��˖�*�ZEA7�P�X�e��"O<)F��5���Ҥ���PG8@�"O����̀�q�)�!�HO�*\�0"O����b�"ݺb+��Y�BL�1"Oz��q�7mD0�8��*mZ$�	"O��z�lJ2w��hȒ霁vN�`�V"O�|@�$�&ԩs�Г,�qZ"OLM��iD�t��8$I�8��1�"O�b�lM�rZ��u��2朠��"O� � A�C���J�` 8,�i�"O�U�X�?�0��@Պ}}2h�"O�a���&]%��!ЮӢ!u P��"OR�IG.ݭ?q�4�-WXI��`�"O�X��x"d-�C/���"ONj�/4T��9X��ȼkvH8�"O��5����ؼ�P+@=5̪|%"O
Mk�bM3�����Ű\��"O��c�ꔒe��Y�bHN�+�m�f"O�y#��T喰�#��8�ƩqT"O���f�W'gX<�s[x��]�g"O2ɹ�]�XL�	��	��b�[�"O�I�U*�u��E�V�Pt���qT"O�����ÿv���#��1{�Vh "O,�xfnʗm��]B4�:q:��cQ"O$ũq��Q4��94)��W�`�P�'o�8��g�@%<�Uj_;)���A�'��X�s�9�>� �r�VT(�'�qA��eڲd��
Xd)2��'�����*0=� ��2`�L��'�F��:Pp�2���Q7@W4D���D�

n�����s�^��#�4D��Ѣ��4u���a�$RZ����s�/D��ӓ��7%WT�z���8 ��yg/D��"w�^:p����6Ξe�)�`'/D��B��Ȃ
�\�W/��$~hPi@O'D����BX�?S�=RG�I�0�0��/D��
�.؝z.��lI9L8`M�4� D� (&e]� �jóFQ I�N*D����� ��r(z�{���Å'D�hX��
j�4tc���8mmHu�h D�<�oV/uۚ�PR'�D^5@e�=D�x���T~�� ��G��@�wG:D����d]M0��%��t�41�n8D����Lw��C�b'�jk�%7D�47��)t�a�KO�^�h�0D����M	�vFP��l�T��șq<D���C�.�yx7�D�*; �b$,9D��Qrh�:\��곇@>.jH��E*7D��k&��o��eR�w1��4D�88���S�,q۴i�y�I�%k4D�� 6���*$�>�#o��ZƙJ�"Orɳ� %��
��X�+V	�2"O���d��6���+���zH	�"O��#Y�B���9�34;��)�"O�Q푆h��B���a���"O��P���^%h�o�Q[h��"O��y �-�.x���#$�B�S"O�Պb��p��u���Oc���aa"Oz4����"���A�g�T�q"Ot�1�N�:S���@&@�@�"��"O�x
ĉ���Ex֪W{v<��"O�"dm�)~)��z���'Vsظ��"O�-�w�I#M�bQ��I
L:�#"OD͉��\�l��7fװ?�T�c"O������twZ�U�>fpz�"O0�U*�Đc409j�"OnQ %��,/�}��D6Z8۳"O�aǈ*v9�L85�� 6"OT8ђ�=Cn$xC�J�����ڐ"OP�3�*M�x����fl9��A��"O�,��И����w���a��@��"OXlX7Ũ�Ȗ��1�0$`�"O*u��$�A�
РP�<I���"On\J殃) >\�� Xx� L3�"O�)`�B:5p�c�3��hY�"OvLϜ.#������#y>��u"O�m�0ń�r��Y�D�d��B�"O��a�H� @�qi�fѫ5�*q"Oc�E����a�f6O4*8!�"O^D��"��S����D�"Wx�4q2"OJ�P�+��ms
��r͌-:�6p٢"O�M�����t��!��* ��<�"O�xÁl:4��ձ"I��y�ذ"O~���J�*��)�e_�+e@���"O���*ľO8�T*�FX_�5(�"O�x���=��v�]*q�x�"O���EIAŪ��2�	���(v"O $�u�v��٠v*Y�6�.0�#"O"H0��]�im���	N�r-r`"O����OQ"�e0�C�Lcڌ��"O�9!%�#!G*�&$zM<Tg"O��at��_����+B�I/��`�"O(�uI�n�⩐Mg*�m�"Ob�@A�$d�U{���$<*���%"O�q�T%^�|L�L�ʚ�?R�؅"O�j��Y/�hT��>� ���"O��sv �q7n]��ǎ�V����"O��1 A�g��f��Sٶж"OD���힡u�ڇņ�e����"O~0��/��M3^ �Hs�\�j"O����(�J%�`�����{�"O���V���3��{u �<cD4�T"Od(����
zȠQ �=Q�d��""O��iB�B�:(�ER.3>�+�"O���_48h����M!0��!"O2m��O� an0t@292�Ĩe"O4�BF��:d�����ިB$��"OL�r�X�x�KF"X+9�P<�"O���%P@5�m0���|���"O<m(G�K��Q4E�+�.��3"O�)�v�A/R9q��AT	+ê]�v"O؅���Y�X%��9t�*GK���"O&���˓�+cڍ����,>AtP`d"Od�P/ӗE�4�!�)��"O� �U��h�M*i3�@7|�I��"O$���
�jv�I��lM�1l�dy�"O(0��'�i��q ��xL���"O��&��:o# ۰�q/�q{5"O��@Rb].`W���q*��">:�"O�ݛv`=:��K��
Y�V"ODP�"O�{�Rh�mf�XYz�"O\�ӑ���W.���؍X���QV"O�e�TjL�v�E�K04���� �'bў�Æ���V4���L/�ʐ�o2D�,"��x�hR�B(X`����[�o�!�ĀyҮ4�r&)zex��&D 3�!���@>���Se��xT��
�DL(�!��7� �zV�K�:6
YԠ�]�!�䂧�p=�Q
�:k<BY��-�!��Y�@���e�Ɠy��<�R��9Ct!�@�~��q0oK��0@�J�:_h!�� ) 9�J�7�^�r��T!�G$��jՂ�%�@3G	��*�!��=Pþ�K���" ��+�C%�!��?Pٮ��QI�y�h&Bv�!�D�s��#���[�V5c��$z�!�䚫EX�d��ɇznB$�I��!��u`pbq�а0i�0{���J�!�$�^6p��G�	[��A拚�!�L.�l�B�%d���j�CS�!�)}E�Dz@�O8ȢW#�}�!�$�{�8H0C�ự�Ғ>�!�o�
U�'� ���iB/7Q½3�"OD�)#�$'P����g[�PPb-�"O"zEK��'��7��5o14���"O�!��z��q�QEP$$��]��"O­(����W�va@�T�t��(��"Ox�0���)��"��C����rB"O�)��cJ;}@�(;���R�Y3R"O�<"�
�8��ǝ�j���2"O�hIgMB��nE{6�_x;\*2"O�d��Ė�5��qǄهg�2�i�"OZh�C��2��ӈ,Ϥ	C�"O`8�@]&f���h ���j�"O�$�["1��
��� V�X9h"O�,�4J������ }Z1"O8��ǻ���cJ�hV���"O�����
W*H�����I�'N��X�c�T1`����!o��[�'�69[0BC�C���(���^�1��'��L�cE<{��,��	��'�j 3�'T�5����>$��mW
��ы�'�.��`�ۯj�#+y&�b�'s��B�X�]�"�3p,�|q�'jx[L�8
@��!HF�vj� 
�'��đ�g5
ʸQ�> _B���'Z�p�.U�c(�%� l�+#�,��'�d��Ҏ]'=zH�J�ɛ���=��'�M��B�11�l��g�I��ܱ
�'�$�[�N1kBQ�P�O�2x	�'J�yf�� ������,]�I��'$���k��Mލ��������'7t�VC�(Ih�z��!wM����'c�x���!��Q��+Mt�����'ƒ@b� ���I�px�e��'�d��&���eF�9��� o50DP�'h�2�� �G���Hע0,���'\V`��n�(QgV�a`*چ&
�TQ
��� b�u&Ң)��)��/R4 l�	"O��r�疧v3� �OR>��"O��x�d��7_@�+��L�m�X�9�*O���`>*t�h#�N_)���'��h9 ��o����U��C���A�',�%�aS/?ƒ�1���:��#�'�5��*�4{/���b�8�~���'�.4a��Z."tv�Hf�]0)��M��'viP�c�1-�B!�"FB�m0�'�&�{!jG(�R�z����}���'��E1��u������%�t�z��'7x�iu.�������m�/� �+���OT��t�)#�jU9nxx$�r��,
���60Θ	ʥ�ǙRɪ�zĈû���Zܟ�'��^c*���uA(|��Ԙu���F�۴0��4*��܂)�Y1ШE�PP�������s�Z*���
4@���a�*C+�OJ�d�֦u�	z��MKCl��C$�P��+�2G�԰�an?����'4��� (o���1"L��g��I�4�+s���zӺ�?��$tr��p�i�	����pnl;�$�O��$�3hv��A�O*���O���ƺ����Má�=Id�f� +��ÀXs��3��S+P���+ C7(MB���O�Gx�C>���TG]�
[��1� #)��l `�8�{��3���I'W?����Q�8{VO^�8�Ő���?3B�������D�+ns��'n�O��D�O��[*�{��F�`��U�=xx�1��Q�\�	����)�?���<�D� �hF�����޴!��7Y�9&��S�?1�'��� ���<-x��:q�ۼR��A�"C�F�����';�';N�2-��'��b��w�ĝ��&)lX�4�B�U�D�X��3]D<u3��y���v�	V�'�xmS���5�L����R��q��Ʒ	P������`�o
*u�|�c���O�cC�'q�&�&eHZI�'�ײ%���`'"5b�@&�0�I؟%����_�4�Y�n��M,L2�C��7a�ZM8
�'�� B©L�HA��0i�9Z(~�m�ԟ�qڴ#,�v�'��6�V:��mџH�I��~'fM<dFD-�b��_����@�pb>��Qd�Oj��O�y�t�322���aJ�i�ޔ��g���CQ�������\� �ٓ��*�HO���C�U�@�-�7m� hx3$۴Os�("#�)F��\�`L�&�yQ�#2B�P#�m$�dH2��AdӀ�l�ȟ��OV��R񨉕$*���� H� ��-8f��O��b>%%����K�~�@���)]gHP�GG3�O��mZ,�M�޴{4@�H@�1�H���b�.Qٴ�T����źi+��'�ӓ\,����Pm�{��L� ͛yP��&jǗ�F�0��@])T (t ;^î�P�lG�
��|�D�O�k,ӭ}f�#Ǡ� tRA
�C�%t4��D�k������|��H�H��[`&����<���5�	/'C�D$.�00X!À��M��dHڟh���M;�ˈ��I�,-J�j��9�p-[Pg�2�~R�'�{��i���F�V�
`��@W�|���Dz�baӰm�L�	3D�[ ���A�T�|��6�
2�5��ٟX"�� d<���I����ܫ���7-�)��I� �K���1�7Z�@�����B
"ѧN��^�.��?�QG��
(�E�4+þ�2)�Bl\�>͂9�1�P�}��ԫ�,�%��5�ө�~�Җ]��� w���~�O�'&-(Q����H�w�F�:���S%x���ڦ��UW?��&X�x�E'E�*M@�� Eј z3�*D��3�W�X8�����u�J��E��C�֯d�,�O��'���M�q�� >  �