MPQ    �Z	    h�  h                                                                                 �L=x���@��$��|�}�=��s_�Ύ��4NѮ@�V^Ӧ5�/�����"�%�V����m�*��Gi�)�<H̤|Yni�؟y�����E[��9�n�uU�K'�u��6A���^h#d��eF&�~Gh�?F^�^��L��h+����t gGhi!�2�3i11ao���(AV�3;u̘A�c��?���L�y���D3�⾁w�������M����LkB��~g�-�Q�Kf:e���F������^3�c��A*T�93?[�A�.��\�-���(D���Ro
��Q��Cnl`�Y�OP����%��ǌ�TV��l?�#�.�[�_������fu8�]E>;���?���b�3cg��\����ܽ��G<��)c0�K�8��D'������AJ�;>Y�V.�ݞ���?�38{t���}��U�d7��,2�[p�~�i1޾\�����qDgD�Pv3��MA�[@��9�j[]-XR�}��w�RH�(�'_"�w��v8��rmq�E����|s�
��Cɀ�H�>#���6Զ�0r�w*�]q^?�H������pZjls�����ׁk�5V����˿O��2���e�3��v9]�����E��aX"tpT�vÛ����z����
��+!Ja�=yQ��x������ tD�H��~m��I�4Յ�'x��zdD>���e�~��T[��l�{�=0���,�=����y��q֯�^V>f+�"B��QM�����S#щ�9o�r+�;퐇u�����]aI��F!�RS&����=n��[�xM�_�6�$�r�'Пs���Q��I�zk1�7>F� �*�)Q)���x�:�a<����pf� _��"� i5������*���f�-I��S3R�[k=ͤ�O�%r���K�"�)d"�!��QC�|Pj���]� ����W��9����"�0H�D7���I t!�2����z�c>׍��Q�-�C#C��ESǸ�Ć�5�V#��5�uEY��D����p��w%�/y$hY_�bS� ��hFjm��<����?�;�ԏ����o�J>}�7���>}�t6����s�e-��م���I��!��X<O�Q�&����|��W�F�]�E��"� 9�_�ֲ�k���ם�O��
�	���U�Rhqwjd�����br�]����*�M�YZ?���+�'[Mg�dR���JoT��-�a-ڿb�T�*�|~�7��I��;^���ue������\-X�V@E�<
��}]��˖�]����xv��O2/�Aa��d�E���>�w�.,R�ܨ��k�l�����m +�6nb�
��QDM��kX���
��:�!�/am�J"�a4�YeW�{��N�,
HU�9�װ���p��q<�3������oƒ��-�E�����S]:���v�n%�W-C�a{�������>�/[�0�9��1u�S���&g���h	�L?ׯg�Hg��I	����|Xr�	G��-��ju ]���y}�N<�����ƭ�S.����q����&��3�?�&��	�«+违���*���z���&��?�z/!�y����|0ݲJg}'��������n�nU&i&��T���2*+Lݪ��2���[��L��2骕ᬤ����J�F�»��<p_�>[l��nq�OtPR����U���_�;o�-�hF���6~�$*�S#�r��el�x�Pt�^�a��7������% ��@j��8�/2;7�#+����џ=�d�����mu��/-Aٗ�[�G:h�jx�ڨ����ԣ&�۟v5=U�]P���L�)"��cL�̆b���P��Ny�B<��q�����Ǚ���~;<	Y��M����O����}���i�>rt���]��{�>��"NF)�(�Z�$ܨ�g�qi�_i<���p6^܉���I�$�q�-�S�%���U���x[����z�,U{����J��f�l>5ĉ�S�m ��h�>�� ����k�ckI�aA|��c���6r״���F![	�XC�wwY~���0��hk��W��>�#.�-?L����"���^�;���Z+��;cY2��?)6�Z��7��C��!���Č�;�t���._Z��M��G�~O�u�1����Ж�@��/�
��{�P�%�����6&F�����w;�Ű�H&C�C�|��#s�\�oA{��L�P浉8���@�J^Bo>�'��L	��X�x�H�V���e�_��ު�t����	��j����`ۼ��ՙuYAN�ou�}FQ��_�,���k(��ᚾc�z�G���G=;R�����9�t(wI�SoߘrD=Nq\���$W�7=�:���ו�ǰ��iS�Z��Mr�`�i+\,���~�l�񊔡�B`��G�P Riv�ZLD�H�lE����uL����ŷ��^I����/*%/�W��da�mÖ+��(���e%�1�8�l�4�+��#��~#y3�͛\b�n׶~*�LY�Y��RC]�V@�杺$�c���F��[��~ e��J�Z�mR��C�E��dcݏ��.���6�#���{��hY�Q��s��
F��8caM1����i;�H��i�L�g��x�**gڃT���n=~\~����2�nf�v��7;�`�s����[�n ��h1�SLgj1p�@)�K:qk�h��p	.�W����_BV�AH�$�7�PO��? ����d�zRϷvM3
5rF�Ω�"��&iK"Cȭ%SJ���i�7��+���	U����)#����@��|di���z�Cd7D'�'��!�("fX.3Ju�D�}/���ʼ�2+����R���Ew`#����f�Z��������A�I�"���7�J�Dv��5��V�W��lN�A��~���`� ��x�c�qM{�8ŉ��g|�����$�$���O�x���5դ]�'�p�&�l��a`׹6M��x*��:��/b�?�I?G/Ը�_��h=\�s����ǡV,%t�@����?~ϒZH���v}�X�����-�5 ��H��DԜ8�#@1�3��JP{�U_~�:_��iO�T�Z�y��k{�4���M|����t��u� ���ej�`��v��UUs���i[6Yt{ b��7���8ci8Ta���\V�2���A� ߚ����q�y�P �r�����w5�g�} �M݉�@q0BF�~+-b�EKA���'�c��������c��JAE�09��[��.�0��<�C���dSo�[�Q-��侎�`��O�ɣ����%	ҵ���Ȥ�V�`����#�	�[���"���a&*̸f;��Z4RB�3>�읂~��Xb�@7G�T)��P���98��l'��腧��<���d��Q �.�-���7���3s�ܕ����gߤ���{��v����l#�
���6�R��l��g�-�1;+M���j���N��]�lm�x_UwM�z��L�z����v�Q��1D�mv���@|�s0�d�#ɛn,����㫾��r#b١X��?F��r`Mًsl�t���5׼�5��E���;O0�}"�N���G[���M���FE���XHwT�nW�VT*�Ȋ���=
�n�ˎ-�J���yL!	u��ϼб�MD���󱫯2�"�o���'�U�z.�+`�einك/琻�&��f0�,+�P[ry�pGqQ�o�9��fS�"��QH����[���{�6��"'��m��Zχ]\���K�R�Ȗ�g=�,[�XL�����f�mD&+��sR��Q:�GI):yk+>��4��h�)L�p�jhƵa2?��e.�pAb_6��r5���x�*{��f��q��3-�vkx���?X�� iF�Y�
K\�E)��!	��C�t�W�Ҷq-X����`W�߫9τ�̝'�Ht>�7�Е�y\&�W�a5�n>�<<� ��OC^`k��Q��I���c#nV������"-�,K��΅���6�k��w��=/4�(t����{� ��Zym5P�凰>�>m���1��KŘ��J�[L�}�=Q���M�����j� �R�����>�:�Ղ����GO����� �v|%�*��Jz����E��H����_-3�������g�8�L���j�A U:a{hl��d�Eө-�}�V�طb˧^3��<tZ���6'�с�b���Q<Tu���<g��W����w.�7$�䊒�N� � u�T�����?�A-��@@�D<e�˫Ӣ.�⨌��\���Yv�bc2���a�#��\J�������,͊ب��K��W�Pm�;�#gkblT��OM��k3n4�E���b��Ȁ��~aO��Y��{��'N<��
�w9�M���+�jqWG?-;���ÛoJ���5�E�Hm�)�:N�ev2@%HO`C���{S���|�{������[?�]9�K�1�S��[&����~�GGޯ��0g���I$�ܔ>mXM4G��w�AJ��}�8�8�-NW���}���Si��M�;��N�āO�3�H�A+	��+�R���[�,Y�銇ه�$�?WS!��.�-�0��P�T}��_�����OA��)t&�H�ϵ0�c�+��.�&���ߋ��*ˑD��v`�'���yXօ�<�]����'_H�������:)�|�%+���R��UKUI�ZX�on��#*���a�����.��`eN�x�tg6T���R;K�O��� ��>�j�!m�*]�7�K���Ѻ��d�*�७9�(kT-�{k�QG�9�%�1�� d�wHͣ �ڼ:=�PߊaL�	��vO����C����+<冉�aB�>�q�"��-�TV����<�j��(ނ���u��}�@X��r/��:N�]W�{ܔ����w+(�|o$m=V���q��i�Ĉ�^^�P �gI��@��w��1�����T�����'��Uv�N��Y�JA�����5?��S�ZՋN���A� ��3��h�kB��I)e)A�c�c��6�j��p�a!VZ���Pxw���Y����bthF��W�Lص��k-:e�9��"[�J^���/��+��Cc��������>�Ԓ$�C���!�a/?�U;�i�K�0�ɚ=���՗�AO��A1�n��KKx@��x/��x�o"����/�|��69�d�&����%;���7(�>=�1�.����u�e'1���^|�*`��En�o��g'l��	�(��F�H��a�e(G��م���Ҧ������&��ۗԩ8�u��p�jX�ثR�/��GѼ��S��y|5���z����FRG��$�E���L�t���.�x��sv=�ε�0�W&�۪�`/�
��.�K��ZF�LM�F`�p�\����9���t�FO����9�TgKRu��U���p�'����r�L[ת������~��ݍ�b�/�a��u�  m>9	������5%.o8��$4>����n��(�y����7�dn��*}�Y����խ�墑3y$�t��B������)�e��i��ZT�(���:EVLxc���i3��VL����({e�Y��UQ�@s�f�F�CW��61�*���&��Y�i.%����$x_s�g�i�[�0=y�}�Z֮2��^n�!+vZt;�T�s�H�Շ1�i*(�Ú$S��1�(�)���K�����چՓ	)����_�uAc�5Բ�P*�?;��<�5u"���
�tF���� ��K]�G�����K����+���	p�2k�#�yh�{�L�g���R
Y 7��e�������(���i� u%���xP��P��I~�j����� m�#�jt�s{�ܾ�i��cئ�\�ٝ���U0�Y ��.���W9j�	�����jx ��r�M��ń�g�i�����?��W��S�V�p�m]JA�p}s�lH���Q�	�-�tӝ܇�?yXbQ�^�DW/p�0����1�\Rغ^���>�%�!���?f��������}EA曎8�!u5��H��D/
r��X��N -�Ń�0��~-�:��mi�
�t�4d֡��4Bp����	�""���u�d��Lj������U�Ysћ��o� ]s&͋��ViS�ae�׃�OHV#R'��A�����-�V�y�,:�f��<8wp�$��IM�.��Br�~Fզ-݆fK��J+�T@<��S���cz=�A`�O9�|[nk�.!�8�cIL�~��D��o�ANQH��9�h`��yO���)Yf%�k�B�`�FV��5�#o�[�먽�@�\��;Tѳu�����3�>'���$���"��0G���)����A��8�
E'$f˅B���7�6���Z.�v�ݔX���\3�I�.+������6F���t$I�^��4A��튧�g�}g����b�*l_�Q�!�gX��dJ]c� �s'ow���ʞ�Z�������,ݡl�m���|�|)f��4Hɶc��44�f�J@Ar�l`�SS?ac>�-)E٦�cliX�賈�����5�R�����Og`��8v.�i`�lve����1<�E(n�X<�T@���3ڡ�@����,�IB=�h��J�DyG�qД7�w�d�+CoD��,����m����b��'.	z��F�:e�}}�
涻� ���0�k�,_����y�q�D}���f��e"x�QC��F����u��ݑ�����v��]����6]W�I���R�^K�+R�=d�][�X����@�A��h� �js��QU�I�udk��l>����`6g)G3��#raMb$�അpt3_q ��6��5�ZB��\*6 �f*��u�3�Ak�����4���ܴ��K��)���!��}C½��~ �Q�S�ܟL��W�,H9�h����HO��7�G���������}>&�{����C��E�{�r�ה���R�#)���A�k �����/��J U�f2�w�*./��-��c�Xĩ �r����m�
傾K��:=ڱ��
����:�%���B}$c����*l�B���;I��[���P�u�=�K�����oOr<�a$K�;\)|��)�̣^�2&E)������_����{��N@��/��ڛ�|�QU���hg�jdq[��d�����SwC˂,��ƂZT�҉�'v��ڑe��x�T���@���=�3��r�e7x��M�c���u[�M�c���z'[-��9@;G<��!���C���J�S�٣}U�v�2e�#a҉���o�\����w\,Hv��jbƗ��w��t�m�lA~��b'�Ԟ0�aM�ktH��O�O�4^�D���Ϸajs;Y[:�{�1�Nwj`
~�d9u��f���Gqr��ƀ�~o<!'�c��E��m�֢:	��vM�%�f�C��u{��m�ښ��%��u'[��9��1k��S�9�&�s��ZBo��9gx��I?{���	X(�>G�����I7�Z��m0�(Nrjo���A|�S�����&`��:���r3<q�\Di	�)�+���J� ��.������?��!�̴�70�N&�)�}]�����<�䲓&�2�J��>$(+�g��i��ڪÜK)0�[��w����-�����������9_����r��&I��C�����U��g�U�o�c�������ͭhk�	b�Q�e�:Cx֗tµi��v��m�������I2�>�Pj1yY�%�m7rX��]�q��w#dw{g��N�c��-w>�g9G��ߚ�Y�����㱣�x�#�=�1�P�k�LA
r�1[��m-��f��;��;�Br�mq��IJQ���:�<��(�?3�A(��}��$Z5rꦵ�U�a]Қ{{��x�K�|�"(�T$Ⱦ㓓�@q�^�i2��9��^R���{EI����'$���B����R���'��ݰG�Uq�6�U1�J�d���'�5�$�S�g����A�t�� �(�Vk�k�޳IDj�Ar!ctF�6���T!Q�ٿ~�w��fY�v��&V�h!>�W�Y1-5��ϔ�",3^�я�o+���cϤ��u���B���Co�o!�'��;�"X��1�d�X���\���OUI�1�;��t@�;�/���
�d��ۏ��7��6T>��8x��;z|�~i��9�����9��/��	~8���+TԢ��U�@��o��''�	ƚ#�n�k_��	be�NS�Ԁ�*Ga�a5_�=�����r�s��u�k�e᠄31��j`�b��a�r�T7@��*z.����גG�{w� T���Et���	+��<=��X����W�����I�%�u��j�uk���3QM�Y�`���\���rv�'}Ρ�{�ï�a���jR����PM��x���˹�f�L�N�ȼL$��M<z���/���͂����m��r��\�6H%���8�\Q4�t��v܁���y)�͛��nMGi*T�Y�ߘ��>���I���$��Ѡw��2����e��dG�xZ_c�d�E��wc������,��:�_XP{ 7Y��Q���s}$0F�	��81��-�Zs���iI���]�x:��gPl3���*=t:�ߵ4Z2Y�un��'���;�h"sة�"�^�dt�$�S°�1�t�)c\K�pbᗅ�!�/	$��>�	_��~A~��-1�Pzd?v�؝��zp��,�
�z�F)��a%�/[K����[�����n���D+l�	��T�%#k9B��o^���#���ye�<7��������(�#��ku�?i�s�ˏ�k���y�M��H]����#<Ӆ�k�������1�w^�������Δ�]�K����W� �Č���З���f �Y=�٘�M�_
���g2K �f���Z*ͥ�~W�.�����*]�z�px�l�/��o��lN��=K�x�,�zv�b�h;�?��/�"����'�L<�\���ؕ�	�G(%�պ���O?�"ƒЃ_�� G}�I�i-��A4C56h#H�weD�����c�ip_�@ׇ�k�~h�^:��0ia*
- ��'@��Ѿ4�n��	'�]B���9u��@X��jB����LU�s����ߣ���� XFcy4Ëc�inra��샦V^�[F��A��E�P׍��y�(`�Q:�s�{w�"�ճ#$M������B�a�~a�V-XQK�'���&��<p���L�o��c5��A{j9�[I0Z.\Bu����ُ���o;G�Qc�(�/`nI6O���+�%���ǝi7>��V�%���#J�[3bܽXT��W��n6;���:%8�3�X]b��¿���~����kGmD�)�}	��@8q{�'_�a���)�2��LK��C�.��������2�3��)�ɩߨ�멤u�����������%��o���t��b�gU� ��KE�:��e|�����]��k�n%w�@�Y�*�@|�w_�������mB�D�w��|�x<�ڑ���xL����a.M���rY���N��?��������<l�[�����2v85'�Э�F(O�Ȫ����ބK���{�r~�lzE�n6XP�T�u���1.��~�wP{�$_��xJ2��yB�+Sx�2��F�D����y�����XX�����'�dz�"��a��e_����ͻ:��L!0��,���zSy3LqG���Shf��G"W:Q>Bj�5<��C���_,c�����&nF�ޝ]R
��W �R?D�F��=߰Z[`x:�����K�cз���s��QpI�I�;k />�����#)B��� ��=ah�h�[[Rp��_�1���5�ƣ�.H�*�V4f3X�ggf3���k�U��u����H��VK�g)�
!��C���-�	��9N�T���pW@��9mU̓�H*�7:��������x,���>(����h|n3�C��3�-��,��F��#�;�dR��=���z�j���+�a��w6�^/��v�NΤ�,m e�	�?,mk�=�}�4��'L�l/�%@cŎM�� �C�d�}��ِ��㌅T����V�����`�j��ư�:��^��}D�O��ӏ�V�|6U����m�;Eĳ<��_��7�6�
�)�`�.�]�����+wUpN�hb%ud������&1��V��]���p�Z�*��:f'l:�ߕ����nTk���:����%���m�7�gz�l��6!u�(�>Ƶ˵�-)�?@6�<��IN���Ё�#�X%vTن2 'Ya�c��N��_���,Á��E����|���m���'�b�+��K�|M�=�k�죻0���yz�r�3�{֔a�Q�Y��{[SN�V�
P�9\����n���yq��.#�ڀ��0ow)����E}����Ǖ:��#vh��%>�
C��{ɞ$ݲ#2���K��$�[�ǀ9�i#1��Sf�&��9ǂ=���xJag3��IZ�܊�RX�G5ק�wi,�������<N�������WŖS�ɩ���\�����7j�3��.w��	���+y�	����b$O逹�7��?͕&!/�r��i�0n̋�b�}�m��������&�h��ň�M/+�IS�\56���ќ�GAE�����������<����C����_��QoY��3ьr���nW��S*U�x��P�o$�}������B���@0#�re=GCx�7�tU��o���عE*/۶��y�&j���� �7�"M��+��D d����[��ϞA�-!����9GK�暛���+q��m����8`�P��=&PP�l5L�*ڻ���um;���"���PB�aq|�x���ʣ����<z�޿��|�����}�N-z�Pr��?�p 4]M7�{��ͳ���ur(� �$#`Q�Nmbq��9i�s����^�@Vu�I�(���]��ZV��V�
:ېi�9btR�K�*Ul����(�J�G ��a 55�Su�ϋ�|��� ������k�L�I_�A��}cO�6#���8 !LV�i� wF�tYφ��ifh��*WP�g����-0� �"ѯ�^͌%x+`(c
������fc�HK�C*��!�5)�;����v���q�����X��O��1����A�@��5/F�ҍ�ϳ�h�6����k6o���Q�S R;X�Н�Z�4'���0c�V���������fi@�`�D�;��oOah'��	�,���:2qD�|e^v��ϛ�����yԁ��ť�M���$u*�=�`�ń��u�%��}�U��
@�/��a�zɦ5����GNLJ��/����t�:���;�I֖=K����W����N�@� �$l�P�<��
MC-�`��.\=�˯d!�B�ס<�Ê{Y���]R:��K"sUaם[��{LQ�Gȗ�;�WO��厍���/;:߂������m4�h�[P�q�%d�8�4��Q�A	o���y��O���n��,*�ӻY�R�cZ�� 5�7�N$m��R2`�m�K��Ee{<��7Z��2$:EL�ccn�c��/���v�&�7�{�6�Y��Q��sXFNVP4CR1{��z���y�/id1���f{xe�g��ő�\=o�0���2Qn�ll��;���sU�9ս��_�<�y��S}��1��)�R_K�O�Rڼ�C	ٟ���$_s�A�o�Ԩk�P�8?���rJXk򛷇�
fe�FD5������dK�S��y������H�+'�C	��>�T#Fl��JĲM�D��^���7u�����W(��0߅*u[��n�܏���ug�PM��t��ָ�#Y-ƅ7��������`�Lٓ8+������_��R�~�yW��>.X��ׄ`�� ������MLNw�zq�g�L��!���u����Ř�	1;���]���psm�l�>?ے'����#Э�S�ᦵ��b�-��:�/&z����g��\H���pX��Ro�%E���?�!��Q+���};r�De^�|ge5��H�e�D�D�T꒑��y��J��Ms~��:0��i�Fe���.��,i48�c�[�ԟ��L�E�gu�L����j�L!��BU�is�����*� S���by�Ɗi�5ma[@N����V��c�&�A��߫0Η̟�yE0�y�N:�w�{�N�vM�؋�Q��Bwqi~|Î-�;LK�a]���C�Y<�Γ���0&c�R�A�\�9Ik[$N.����8��T!����o�l�Q~���/��`I�BO<��_n%�Cl��nn�VV9Y3+��#%Z~[n����|�R����F�;�(�����23�>�!i�Zx��y���QǓG(G)���7��8L'����x��-&H�����n.�h8݊�*�n3$��dH[��]���<���(�ǀ��j���qު�g�#~S�]K�g�b;b�`
��G_4Wk���މ]�jO�iww^����ˊ�����6��l�mݴ��rY |ߪ"�]�쭈�*���<k���r����I)�?�F��a���l_��i�]�md�5
����OQ(��}ޟV�b3��MK���E^��X�4T�(�ÇP&�z��	����0��|$J�;�y=���1y��ٱa�D����G����NP����'��zPWV�|de��	��Cӻuv�o�0�u�,O{��:�yN6�q�Y<��=Af >"�#�Q9�~���ܧ?����U�Hʘ��
�a�?�+�]M5����ZR�逎aL�=Z�#[;�)�K��w�w^�J<��s�e�Q��,I�L�k��b>2���1�)=m��{���)va����!+p��_�;�l�55�R!׉S�*��DfN���xo3�@�k)�*����$�j�K�i )�F�!zz�Cxu�h-�҇��I�(�L�W�%-9 �K���H��7u���F�w�h�f��>C
��q[�IuMCx6��%���8���L#���^�a{�[�Z������\�w���/e�3�N�� @��ӿm�C�x:��O5��'��@��	!�����}Z���⨌�W���\,�q�A�Q��E}&��.˂�/(�x(O(�סx�q�|������7�nE_�
��4�_>~���N��DPɝ�aػvBn���pU�h]��d'�F��{�΢��IVI�8��9;|Z�����8'���PQP�&'�T�.����Nw��@�h�{75wu��f��QbuQ������*-�q�@1��<v<���:�3 �I`9�3�v�Ė2�yfaȵ�m�������*,>�T� x�����(�/m�.d4�cb�ǯ�fޟM��k�� ��1w����͚}�6�a�O_YQ��{6�pN�bd
���9�b��n�\��q��� <�{7�o�/�͙�nEx^��:�h:	Yv�\q%���CwXJ{���M�A��?H�+aG[p�9)�1a�sSA�a&S�v�ԛC8��ӱ�g�EIu����GXު3Gp����%I�Ir�iĪN�t��x.2zS��\1���1Ē'f3�"�$�	y�+T˸��>���9��{�2��}?���!Jf!�u8#0Ij�6��}����m�`��Z��&վ��@�H����+8��� ��H����N����v�o���6��.V��$t_Yi�*�	�&_���L����IU:�K��olC�T��	�=�=�˿�^<e�s�x��tx��M�|��᛹�oRۑ���1jg�Z���7(.��*�2�dm|`�6-g���1-�#����G��M�V���FI1��z?����ۋO=���PЍ�L�j»����8���m�����:~�B�hmqw��� zǅz���v�<�^���`����FCO}�r�f,r`J����N]��
{m����#(ܢ3$~!��	Zhq�F�i({���i^�p�iI�u�����?�n�������D@��Q��0ZUg���@�JrJ��ػf5�?#SP���d��� �����mks�Iz�1Ah��c*�6^���A��!G��8w��Y�5���h�c�W��]����-+po�J!�"�S�^-����+;v�cE��ū+����ԣYC��_!'���;m����Oʚ8�������O˜�1��ļ(P@rcL/�ڽ�@�����������6��0嗰0.o�;����,��/̂�Bu�_&'�۝�������s桞������6^#o��'�?m	�ގ�d�?�/�e�������[������콗U�(d�B�u�K�[�Ƅ雗��!pј	��W���
��O�<zd�ʩ�YG�<��v+�F�t|�V�߄7�=�ӵ����W7�x�	�j�[Y����$�+�?�F�wM� �`�E�\���jv��]�(��4��ew!�m%R�0ʁFT���)�X���-��L̝8�rzC��ї������/��ĂC�4���m���6��ìB%�C�8��~4O�O���%�*�fy&~�ȕ�n�W$*Ns�Y��Y��L �B>d�R�e$��-���(	�S�evm���VZ���M�Eǖ;cI8��u�'M���� {��Y��PQ��s3 �F�+�#�1v���� ,�4��i��S�hx�|g����,�=j���kQ�2χ�nҤ��G�;d��s�V��X���Zh��Ԗ�S8z�1�l�)b�K�NW,s�W��	.����?_.�mA���#ƫP��?�mv���f÷�
�
!pUF_����2��KD���qa���d��e�+�"	�*���P#!��,F~��.>���Y�70�z�GO��N(�Q��]u����is�a���z!��s��>�g��#�>M�Ҽn�
`�z�~�4�ZA�
�����
����˹y�'WJ�:���5�_��) i�B�O�yM�\<�uSg�mƺ�3i��҆�v-F�䇕�!ހ]Npn�lY�O�M�%���o�����.�����Kb"��5_D/��Y�K{�ɂ��\é��K/Ǎ��%�T��J�?wG��F?;�5K�}��ț�iӷ��5l��H�s9D@_�c&��p|�6�D��PZ~�qy:�Оi��]����e��ק4��e�6E���?��:�u��	��j��̦�u_U�:3sbF$�Ul�ŢN N�/�����i���aִ��\��V�o@|�EA�E���D�y4�@��%�)��w!��AM�ݰ�BFB2��~��N-NFK��Ã��u�%����c��% �c��A�n�9~�d[�r.�b��4����n�U��o���Q����P�`$��Ow�u��0�%����S��'�VTA)�t6# ��[�����/�M*��$�;�����.3k3�DK����`��t���BHG��)�b��#�8'��'�j��q��(�*�>�=.��^��Z�3_oǕ�/����+zgܠ��F��
C]�凵���]�X��g_v�|{������2�:�G]4���d?ew�׆���6���m�ӽ�)e�mx�܀mLH|:�H�P�M�����g�ٶ���r�L�D�?r{��^C���Z�l��g�DAWרr$5]s<��8Ox�%�i1�޺�����̫(����'�E��<X	ثTQ��B�¡4#��m㜻������Jh��y8��/:Ϩ���|�D����_�ů�b�eK��p�'?;�z�ֶ�P�eUl򃛢ɻ�O8��0�*,p��<Eyirq=G*f?EH"IHQ4"/�W����y�	�2"N`��5a���l��m�]H�\�5fR���|�4=�1�[i��t���Yܹ���s>�bQ�YII�kx�>mn��1_2)8Nc���VT5ia��	�Qp�5_"��$�5�����~�*gd�fi]��3���kd.rͫ�1��;��I�KH��)러!��zCS�S����"l�D�X�]�W��u9;թ̉��H�Y�7���P ��ͯð�!��>^9��m�$�CJM�Lji�ȼk��x�#Z�8xl���56�j�௓�� �W��w�р/ i��8���]X :[F��m��!�s����b�����[ ń`�P�8��}��B��j�;���s�ٌz���%� ���&�� �s,�O�f����N1|)0�]n,��B�E�J��u_�,����I�_z�$6��Q��-�>U���hX9�d��\ӕ�ұ�>���un�ڶ�t%gZ%�B���'"#�����A��Ta�Ш�S��l�[���c.�7����~�z�l��u�j��o��+��-_ys@,��<і���y�N]5��`�%v���26�Ka�{��ȟ���5���m,�� ��2�7���í�m���habX�c���M|Jk�E�1S� eL�(vg��C;a�m-Y�~{?N(��
O�}9���wtP�]�që>-�V�o�f��4�_EsP��
::frv�P�%4meCR��{?o�������솽�[+w�90�1�g�S/&����o��3��.9g���I�y�܀��X�g�G�g���?xZ��$#$�\N�)���jVu�SUp���&���x��p3m�U�Ĕ	��g+/��������o��vkH���?C�
!e�״�&�0$(q5�}.�����헻N!�/ &�4ջۨ���M+s2H��,Ƞ�Ǣ�\���x4�1;M��.J	��q;^�����n�_���+�A��h$�̞�>h]U���F�Qo� 	�E�$
B��Wh˚�����es�x��Xt��j�w����;�!�l(֮�>pj@o�I<7�O�al�&?rd�,���k���-HF+��h�G3����aA��cv�m����=\zuP���LR�*�b>i�S��kګ��Ӡ�uO�BCa�qr��Z�~�@q��ER<p�o��!e��\��C}���0�r̠��r�]C��{H���f3M�(�D-$�͓�fRq��(i����ʢ^��ȯI���8�ӟ�i��Ur �����N�݁�!Ubߖ�fw�J-mP��5U5+��S+N��:m�E�U ����g24k.��I�9A�śc.�6��(��?!B���Iw��Y���h�&W�ȵ*jR-&	�ϥٔ"G^H#��h+�c����F|��R���C�:�!B:+�@;H�7�l�5�����Y��"O�v�1
��7]0@M'3/�}������#����hbl6����0�	�>;��T�O�m�*�����C������z}�������T�����1�!o`�'X�O	����ܫ��"�e�%E��1$;$Ғ�{
��f���f$�{u`k�V�D��.ѳ����A���'��-�z�X��J=GMp�1G��+ٶt�g�?߿�=U|���`�W� ���;q�v׏��o�^��x�My4B`��]\��%�éxX¡2�G�@���@�Rp�؁A�����O�H�LGu��MA;��s�� ��n/񒪂��Ѿ�\m*������?%���8ƴ4�pm��� �E�y��X����n�P*�2IY՘T�_q���בm�D$���������eq�~X�Z@�k�h�EB��c$�|�U�H����
D�i��{Q��Yt�Q
Q}s�F��j$�1q�w�0����Ii�����y�x���g���Ǆi=ew����2�Tn�e�b,_;?d�s�E�����U��/��S�P1��)���K�mU�&����	�<�O�Z_�4�A�}�Ԟ@P�w?'s㝨��aR��=J�
ܚ�Fz���Q;b./KITO�,���������'+��	ܗk�#�8��ga��������v��7�J��v��(i�U�u��$�d�L��5����͹��댄}#�oh�m��ǔ�o�Os��Ȉ�ى�N�~��E1��}}�t)W����;�P�/�VO� D]}�M��Y�pU�gC�麗�������_ÿ���\0]���pi��l��_��C���L�U�	�{�+.�b�b�0��/܈R���ɝj\>���&�	��)%{�֝���?�	��M��Pp}1#W��4���-�5��HաmD������� g������s�~�:fJi��q9� 3���B�4.�s���~��{�@u���i�(js�����Uy�)s=�㫐 �`�� I���&���i��;aQI��7V�
A��1�aC�B	yO��&�=���w\��Մ��M�R�B��a~�1�-�pbK�5:�6@������S��cf�4A̠[9�
[�>�.#c�ϧ���x���olGQ�ѣ�%�`�XLO�����c�%�/�Ǯ��omVoI!��#�/[�/�)͙�H{���;@ u᳞���3�j�<i��o�>�ޜG��r)!�K�-ŗ8��'W^����#�I�]�����.4��݀J��5F�3�fT���Z�ԡ����"�����%�`B8:�� ���Y���S%�gf{��A�(��=Dw�V�u�]ϳ��_��wZʊ
s˵�g Ә�X}�mԼ�h_,|�o��k��"xY� ����E��6Ur*��?ō?������8lU&%�����5�hf���mO����$�����Xp�'�a�E�0�XL?T������OY���o��%�T�^J�2y3n<N��co_���Du}�:��YE�)����z�'���z� ;��\�e��F�v!�����=0���,�\���y��q��+��q#fz�f"�3Q/�{ﲳ}���n�$���s��]
��^��a�#]C���h��Rp�Ǝ�Ɯ=P�[�����E���}T��s��SQ�NI��JkS�>���̬�)3O�1�ia�a�.f��p�_]�@����5��p�?�*"Rf�����3t"Ok��m�Fʠ��� �iK͆)�!p�gC.���[ҽ��?[埸nWq��9V9p�mLH�0�7�Pܕ���-�}]�)�>y��g���X�C��w����ô:�Wp�#�{S�u�WVfͪ�x٪����R~�wG�q/����]��D&� �|�Y�m<5��n6���ڝ��vS��'���hs��}�9됇t'��(�.D�٧u	�G�r���<�aᨂ�0��nP'O�	�M�6�4�|����8G��7�E��O���_��Z�gb��z�r��*��,*��h��UA�shS�d݀R�P�����?����p��/FZ�H��iQ'}G�ƐK�\U7T�	�ЃhϿā��e[�^~7��ˊ9�ƇfuG@����Q�f��-���@'ɪ<,��z?B�i��?�ɣ�Tsv��2�~	a�a�#Et�HC7�X�,4d�����r�C�^�Gm�pw�8�b_���d�M� �kz�9�l��������q񃬪a֫#YG��{�4�Nc�8
�jK9�Н�Қ��NOq�Բ�y�1�(o(�'��.�Enb	��[�:��ov�dc%��C-F�{ze݃����ٵ��9h[�~T9Kn1WJiS�@&�hi�
��.O'����gdK1I�c����5X�D�G����H�\�'������RN����n�J��0S��Tc��D��H�3(T�Ȅs	ow+
g�6;�3���qtZ�H�2?���!����k5?0��΢}�O�������X���A&�v�655�e+��P�-X��fe��b	r��L��᎟�%=֬�x�dc����_���w1�\ڌ��r�*�y"eUR��A!1o5���ʤ��?aέ��u~�Ԧ�e-�x��.t.� ��a��E��Z��G]®*�j�<��7�A��I���Al�dc�������Os�-�7���bG\�<�̜��|Y�ޑ}�Hy���"=�'�P�/VL�K��a�n�$��@��r	8��@B�y�qm�a�7#���ĩ.3�<롊�o֧-Y{|*p}�ӯ��#r�mw��K\]���{#��7n���q(��$4ۓ� q��iꌋ�٣^>�'"nI�o����!��#�{�����l����U]7����OJ����5��JS�/�u�e��� ����´:k�UvI���A^�\c�et6�*��w��!=�̿zs�ww<�Y wX�d<h�	�WD���o�-!�@� ��"��^c~��S)+�q�c�	���� ����Y�\C[��!]���;#F`r>�Ф���Gїi�OAp;1%$#Ĳ�\@(�/�x�vC���G5�#��6������l�;	c���o��%v��]��%%��S��g�nf�i��1���,��o`�'UV	2���Z�ˀ=���e/����� ����Mc%�������c�_9�u�ƈQ9]�����VcQ��y�M1��b̾��-z�_ݩ�[nG_}���m�F��t
^�u��Y=�Ds��<W�{W��u���0���V�$oMh�`�sO\N5������ᣡ�mZ��!�{�0RN?�<f�Z�Α�cw:L�l^�((#�6m�����S�/Lo���as���m�E��쥅�"�t%5�8��4x��r���`[yy!ߛ~�<n9�*��Y�k�t��������$��@��J�π�^$el���b�Z��6��$E���c� 1�����]���d�p�{�Y5 Q��js�[<F��E01l�ϋge���Li��\�I3�x���g<�b�bD=`v �!�2E�{nG��0;��sU�Վ���P�䊉�S���1�y)���K\���@1ڍ}P	8E���u_��lA�4��� Pqa?b�d�CP�\�巘�
��F����7�=ÀK��ӭ������J�YZ�+X�N	�$�}�#�x�����T����ѣn7�w}'���%>(D���u,���_���-����H*[�4h��g�#
����� X��0{�
�����-�#�YY�΀����`g�o�8W :���S�k�G�ѫ I���uvM���kw�g��R-d����l\�Ú�����]Q�pdԞl�p��f�ؒ���G���`�f�RbX;��+�k/7@k���ɸd;\�}�����%TP�0�?-촒�z'�k�}������p�-��5���H��}D�3���y���9�,e��w�x~T�d:|�i��vNL��v���4�ȍ�� >�I'����u��C�W0j.Y��U��KsXS�˴���� DB}��Os�iڈa��:�cVJ�u��&A��߼�ϗ��	yjY�����ߦ�w��$��?M�Go�b��B�`�~͘g-D�?Kc���q�[o1��c4����c!�A���9t�[[��J.Hp�j�g��>��o'��Q�]���`�HIO�lW�0��%����	?T*)�V�q���`#���[{3�Ċ�C��ڗ�;�����,$  3`�yNń�+��j���b��GY�)<�\����8�~�'KcŅIx��ۤ����J�.O�L��V���3�}��5�ި�s�����5=��m�ۙ[�H�[�-��Z��N�
g����	����������>�� ]j���Z�wo�M�E]�)6�cU��s�t��Dm�U�c��|�V��H��=�����͍��qP,rŁ��:�B?(�$�����-;�lЩ�������5�~�����O.��������7"��>N��ğ�X��E/��X���T�øl�j�^�c�n��nǎ�I�J���y.{����yȱ�HQD�gO��3������I���'��z����͈�eK��Q���&$��T70���,&�̛�9Gy��q3���[�,f�/�"I�Q*�d�s~�p.��?�����8����c��|k]>v���=R++Ў���=�2H[�7ؓ���H��Oh,M��s�G�Q��:I�k.�>���g=).p�ǌ!�ʬ�a����G5�pc�_�6!�=��5��Bך5*��Nf�P$Sm�3OÊkچ��H���{V�K�.�)!�o!�O�C	�##x�X�s:�͟0W,��9q���tKH�'�7&#���3���	�yi���>���������C�����S��̥���V#Іn'���B��V`S�Q���Mamw�6�/�dD�J��t �	��Lsm׏f�i�r�`I�X�A�@s�z[��lvU��>}+��������������y����� Ɯ���Ra��i��O9�����:�|���@&�YK�E0bƽ��_O��"��ó�?�����VUܨ�hN�7d8�(�� ��ǩ����W��YZ[�;���'؋#߁`��w5TW���^b[�����B͕Y�7Fe'���Ƣu�5K���;ˡ(�-��@"Z<����5%���w����C�Ĥ5v@F�2l1�a�gj�~
A����4�,����ӗ�'����m�A�E)�b�ZW���9Mr�YkUq���&VV�)?ތ�g1ra�	BY¡�{ǅ�N�G1
�^Q9�7b�-�2��`�q�o�'��oc5z�j�JEi���K�":�QvԘx%*�pC�{����@���&�<��[���9f&�1�L�SҒ�&� ��)ׯ�Cg��I�m��v//XoAG!xy��'2�}��Z�Z��N��'��{äS˖ӵ���͢�ģ�3��d:	�Z�+�cf�q���:��l�h���?�$�!�g]��c�0���}d0����C�q0��&&��ձ���0-+��ȣ:��%d��-,��g]��	d� ����g��V��b�_jeT[l�w��^,M�����`U�>
�<v�o��$�Z�⭁�"�P(
��e��4x���t���~l~���չ1 ��"�ޮe��j8����79�Q�m��\��d��P���eϊn-~����G��Ú��֗�'�Y���#$b�<�=��zP���L�{��uޙ��6�a�L�M__��Q By�!qh
=hǶ���IAt<fsѸJ��hu���}����?r�/��DO]9�{��C�r����!(��4$�%ɓ:��q&��i�Q��0)^yI$�I���aJ�p�Ё>�i�Cy���N��ݷ~yUX���F�J��)�*5!�`S������{?� �7#�W�k�C�I�cCA�6�c���6~��c�!8�o��@�w2��Y;���[hh�W<���`��-���[��"��z^~��2�+�Fc�rD�|}L��5�Դ�C8�!x�!?;�������k�+������7�O���1@u��-&�@q/2�w�� �EP�����ދ�6�*���P��;D��Aa� {^�S%�U��,�~�pr�Il��R�������'n�o���'��	M���g����0Ce�T�ݻG���;�R�@�O��+۹&��"u�#��L����=�4���ah����뛽� z�z5�Z����G�͖��ު�a_�t�Ta�P��5�=�-v��8vWH���:�j�3�������j����M���`�:}\��˛kv���͡(:���*Z���tR���7�����׉�q�~L=���/��CFT̒�{�&/�kv�t��!;-m ����Wx�]��%С�8��U4`�	�-�"�{��y���YL�nt�C*�Y�^~���ӯs����Q[$�������Y�:�$�egG2��Z��e��dE8Lc��U�˨J��m 6�{�E�YP��Q NdsĹgF:�3���1gB���:r�e��i�����:x��rgw����V=[�h�|��2 �gn#HOXU;��QsA���)�k�KƷ�岧Si�1-�o)xP�K7�{~�(�D	�ɧ:�__��A�Ԕ�}PLk'?�����<�W2��(�
RP{F�}��<QxK�ԋ�b���-X��U+��	Ҹ�m#��4������;���,yk7a�B�-�l��(��^�u��$�Z���r-���FE�ͯNS�B�F#E2[��&;��u���ŀ���D��>#�4�λ	q�Rd��j��W[��k�/�N��L(� �Tc� ��M�H��f�_g��кڷ��>���#��uLE��4)]�z�p_��lj0��~F������Z�ӿGV��H�b�t�&��/���|ca��~\4b����O�>P.%���z��?���w�Ά�s}'T؛��l�ht75=��H�]jDQ:��@�9����X˫R�~�L�:��i�=�Ѧ߿���(�c4$���,������zu��
��j�G��3h�Uow�s�s���Uz ?�@\Ӌ
�#i�9+aG�̃���V���M��A����֐����y��������w�u�պ�rM����Bc�j~��-�%�K>�W��
���^�����6.~c��(Ae�9�^Y[���.���������f=Zo�C�Q�k���`�X�O(xF��(�%曾�d��YYV��{��#��`[Z���_h��>}Y�5H�;�Wn����\3;i��`���t�e<���t&Gf/)Wԕ�#h%8���'�����+|�<��5�n�.j���v�B��3������e�<B���a�3��V
���ޖ�W���L�I�g(N�d��|�3����6��S�]}��Uw�w�a� �W7�H��bL�Njb��mIs��^�(|K�<�F��X�J�g������Wr`LE�5��?�����}J�H�lKMd����Y]m5.�����3O�������C�N-����P�3�E�Q{X���Tb6�sp��%���/��k�Y���iJ9��y)������٢��ͩ#Dk�m��"��C[_iM���4'PwLz<j���Դe�z4�,M�a�7S6�0�	�,�`=�my�y�R'q�L�6%Ff���"��Q%b��hR��+�ÉZʼ�+���M�-�4k]9!��	R�����=F�A[���7FA���J�/��"so(aQ��I�zFk	w�>aS���))�p���[a��7��{p>�_���ح�5��0����*���f����L3*�vkc��|q'������7Ky��)<k=!f,%C�dDT
���w^5�n�W瘨9�a5����Hq>�7a��!m��jb��u)R9->����]e!���C��	��������D#�������M��ǆ��h��%�Hd�w��/Q�1��:4 �!��_Wmr
��d�����8�#��{�����G9��3}��$�}���Ly^��������=�e�t���ׂ��d��O�������`�|�����X+�{E�u��0S_��2���f��<��s������'�Uw�?hI�d�����N��:��5�fˤƲ�%��Z�K쉈�Z'3�>�<PW���T�~��9|��:�,?וT~�7�������ƽ�u=K���^U�܈;-0P&@_�<�eh��*Z��4)�5"���Hv{�2a������m��Df�O��,*����#Y��b��@m�2{�9[b�v���j}M��k07���v4��<��9��"؃a��Y=��{���N���
 r�9�b׈GD�H�q�s�r�����o�̠�DEd���^v:k<v���%���C�4{��ݹs0���엒�[\�9�eH1Mo�S��&?���@.8$�"�?�g���I�l���XJ^_G\00�~��0����VU{N	r�d4��l(SZp��F��� s��\�3��d�	e^P+������e�i��g�r��^Y?t��!�R,�a��0�!�"a}�0�����̨��F�q&AW��,H��`��+$~�cȠ���m�v�3�4�H����"�*���v��:_�N����O���J�(����PU����7�co��Z�@ď�uo��fR�+�(J��eDf-x�7�t�Q��9��*9��Ř��&+��ej�&��
�7��2�"��w&�dY����Z�ŉ�-nإ� G���B��ֲ�I��(l���z�w(=-��P�QLc�d��Aߙ�Q��m��(��&��B�qcv4k�L�q%�doA<�dD�%$ȧ�����q}�!�A rLq��]�]�%�{ه����*(��B$�f���LiqA�i��[��^��H]5SI���I��+���Y±q�������R�	USGt�w�vJ^�'�Dd5��"S�T��E���2 ܚ]�xk_Q�I�(�AT�Cc�516J�,�=�!3��0.Xw�M�YV���ghC/TWw ����,-�϶��"x"|^����0�+��>c1�V�.������\�C���!�l��X ;���������Et���O�Õ1[��Ĩ��@�2�/m����0����G~��P6����n3��*;� 3���J��ƕK�3�G�1�뜫$�捳��gH��"^�o�'���	h�F�P����kfee�ݶ�L(�÷�[ӫ��G۔��կ�u1V�G%d�U����$��j��C�v8��;P�z�zЩ���G>��bZl�|Rqt �p�+.}�p�=&6���T�W������]����SZ��p.�2�6MJ/�`{!�\t��V����S?��&d�Ѧb��RA��2\���D�ع��gL��4��U÷~� �v-=/�\�/�¾<�m�*l��){Ø�%kV�8�,+4�懣��i��O,y��4�}n��*�1�Y�q��*V�.uʑ�ƒ$x�����̏��H�S�eb%Vi}�Zq3����E�d�c����y��c.���z��{�Yk�Q{�is�7#Fu4_;�<1b���A.� P?i����?�x\��g�%�Ř��=V���
!2�nn>i�әn;��s|�u����Fм�@�MS$��1H��)���K��Cտ�à�	�ʧ`��_�|A ��p�P'�K?�B��yI�R�x�N�
�zF�_���a^�L�K�Dx�������!��K+ι�	-��s�9#�X��s��T���,�n�7�]h���|(�<�ub1��U����M��f�`@��*U���#��2�>����u���&�7��Ӻ���O�;��������e�9W��&7���P���> Հ�;��MS���a7gT3��Ȧ����ۥb5�P#`��]�t�pZyl����9�������Ӛ�[���b���!/���7F���{\���ط���y�%L�k�u� ?���26$Ρ�}�˛�\�ӣG�5��@H��2D������]��"lЫ-�W~�* :7�i喖,�Q^��C�64�e氢<������L�;u���z~j�V�NNfU� s��B�A}�1ѣ : ��*J�ņti�a�ƪ��J}V����ghA�mZ�r�1�s�y���������w��U-M�1�^B��~Ǡ-:��Kc�����"���P��}dc�8�A��9j4[km�.�#&꠾�������[o�	Q�'��`��3Oc���f�G%�yǿi#��eV�!�b;#l`1[�Ǘ��e
�9.,̐�;q3�2MaM�3���'��aC��`�z�p[G��)r���i�8��r'�ۯ��4�I�nr�)�.��������yj3K��kA��w����2Sj�N�5�Ѩ$�n3��Pv�*�7�D\gw�c	��ň���v�$?�&�]����P7w%��ʻb R��Y�d�)G�	��m��YXA|��c�<d��s�o��ߜ�}���6�r�6��0A?ް��J&��c�]l���L�ה�m5�	�����O���U@��&nm��; ��`�����EekX�g�T����.ʜ�����Y��F`��r�J�բy$��Mi�ϔ���*>D������
� �����X'� �z�>��A�eAj̓^��x��7�0�>�,�4��(�Yyթq)>.��of+�:"��Q b
��Q���$�u;�q��H���o+�2#]4��yR������=��[�ׇ�r!��~��Et �s*)~Q��I��k��>YG(��U()$�B�@�^a
ج�=�pM�_���s�5��:�Pl*S�4f��I�23ekP_���>�����1�=K4R�)WDS!�(�C��4��Ҏf�0A����W�Ł9�%4�u�HLuA7�'U��ƃ��6�/���X>�5n������C6�p�����\P�hS#F�� ��Ȏ ���̐㪇�L�C��wX�/��L����?� �Y�2��m��_���X���ch� l�p"��"$��}a교x?H��QG�_���&rѸ_����]L��"ϱ_|�O�1~�����m|����ɑ�����Ef�[��_&?�������ȳ��u����U*hD�Ad�,uӁ���U�3<�U<�`�Z������'�tZ��_���
�TMi�����u���[y�O.�7��>�j,�����u��e�`C��	�-��|@��<=@��PL��`�����z��v�<�2��Ra�Ӗ�4���y���jP�,�f�g^O�#4 �/d�m�C��iYbD�[���Mh��k�������@�#P�ݞ9a'&�Y�D{}�XN�>
��9�e������	q/����"roك�͠��E_X���:&�v
a�% �,C��G{+Lu�T}���0}��n[VM9�ā1ȱ�S��&zpl�ۢ�����g���I���l*&X%��G������.���N/>����yT�SA=a�%��þ)�Y�X3YU��	���+�i���7��#�bOy�Y�,?/,!�]�� D0�_�]Z�}�Q%���	�'\���&\Mtէ��;��+_���������ȝ��_f�����Lv����]���5������_ X�ѵ�����T��o�*5U#�`�2��oF2!�����&��w��W���e�2�x��Yt?�������*�D�'��ػ���?tjn^�5D7�T�z�ђ�wd�.C�},�� Ŋ-�m�ހIGmH��^1��aT�O�ţ��۲n�=��`P�TL��ͻN-d���s�W4�k^�a� B��q^H����,�K��6<\v� eI��[MuF}�xO�6�r���]/��{�s߳�C�l�(��$E�E����q\��i��:�6>^�a��yI�֜�Z���'�tс����I�ă���1UN���Ҕ:J8b�_^�53�S�AA�&Σ�>� �T����k�I�A�'icq�6����H8�!.JJ��;w��Yq�Y�~_hrFW�����@�-�]���"3f^�O%O�+���cl��Ų�+��݀�j��C���!����;��#��ʡ�;�����z4(Ori1vw�#o�@�v�/�VÍG׷��X
�T56���m�u�Y;�aϝ�D5�岬	���bam�f�S�J�Ȉo��W�n5oq�l'D�B	�9��r\����e Dݱ���?T�~=�vн�'��o�%�ų�B˱��V��5���ɾ/o�Q�ξvF~zk8>��N�Gpν����ejt{!��t߫��=�^ĵ���W�MV�������V�ra��m�(M�¿`v(�\_Z)��9��<��3[ìB;�,�xR�郁-.�w�5���#���L3Bȹ�{��<���q��/]�B��Xp�W�rmͪ�}����%+�8���4N&��Ձ��y��{�ffn�0*UqY������6��RN��[�$�߲�t��8��Z��e]#V�:�Z,���D�E.�Hc���A%�.y;����k{=�Y�`�Q��{sz�nF���f�1]J�ϜAl���.iV����x7:�g�i�3s$=Q3��2I2vx�nY��N�;�ss�B��_E@�A��e�S�!F1c	�)n�OK�(�~O��^b�	�G��B�_��
A;�ԊjP�?�`�vM������
ȅ�F�af�u��A�K5՘��'-��#��j��+��	H�&�n2#h���S����ᬂ�⃅7�Ypx@��bXr(Շ�A�*u���P��(���!\�{�ͥ{����P#�t��ٷ�񻒔A]�;��4���u����!�1b2���u�`EW�&�4�`A�B�B �̉�vk�M�?�\�jg��7����'u����+k�H�]"��pU[�l ����)���{�ukq��sb)i���/H&v��Hu�	�\*}oؒEVǴ %���py ?>S���Èμd�}��fTT��:5sB�H���D������&!#�����?o~),:�l�i��������^�4�$�}��������u���Aj_�ĦiTLUe�s��«|�Y�l 5�����@�i+�:a=�ԃ���V����n�A�G ��貗.\Jy��Nֈp3�wH�b��AM�֯�sX$B�o�~�	-�Z K�\��"U��,���SI���jcR��A8��9�)Y[F�.�c��;�����R�oX�Q �9�S?`k� O�� �n�%܇�/�[�V۩��#G[r[�����u�4����R;,/xM��#:3�A�������}�[T�s�0G�S|)�p���c8n�'�G3��%����]n��.�?��l<��u�3��ѕ�{���Ĥ�Q�V�iٵ�L`����ӈ��W��?Y�g�,�� ���)��yvW�aN+];��K�1w�|��v�m�f���(�D�D�m�n�T�|y�����Ɏ�\�x(�^%��"ڪr�A��+}�?9�c���~{�lA�S苟��ϙ�5d�����O?#�����A9��Djk�o^b�	��E �rX�[�T�h��m��q���u�!	��@6EJo!�yX,�A�OV��̠DaU���$q�E�z��\���-'�cz�3���se�y҃�\���RQ�Y�0��u,7)��X�y� �q�����X�ff�"P��Q���qA���na�Id�ɝ��_]���]/�-��hbR\���;=<��[]�W����^�@*�^�'s�I�Q-2rI|��k���>�Mq�8#�)��ǝ���O�a%�)��h>p��_I
<��F5�:a׫7*6f��āD3�e^k�{eͲ����6܌�K��)r=�!\EC����8~�)u<+#��$4>W]?9�	���J�H'��7�Y�W@�龜�����Ȉ>���S��k��Cq�S�港ԏ�Í�#O���+�C��}������",�>ʔw���/���g2��0� b� m�m�_"�Z���q%8ډ��D�뵻���_Xz}�?�s��J��������3>��g�*�M�U�#��Z �OJ�N9d�a|x�W���E�
H�E�z���_`t�S	O��V'��<���yh�T�U�|lh?�dI���<xE�p+~�+�}�Z����KZ,ϵ�~�T'�v߲�s��1_T�s��`��Gb���J�`7Ws��%�����u3���;H�R�|-f�@u�<�:֫f����_�+C{�UT]v���2=	qa�9w���4�%��8X, R4�B���^�Q���m�toV��b����M��k�"-�X�'� ���Z����aB�Y3Ƅ{X8�NOLS
V��9�,�>t���U�qJ�T�����~�o[j�;i?EZ�f�\�:�Ov%�(%��,C��J{f.���x�ҍb�Mk�[���9�CC1C�ScH"&�]@�v7C/�����gP�IL����#X ��G� :�������k�˖�NJ�^�ZT\`S|@�����Ⱦ|�Ĵ7C37�4��	[�2+v�"�}��[+�]�{����?���!��W�0k��s�}5����2��/w�(2&wcn�"���+��|��F���"ɜ#��^)]� ��zqF�L�֘�,��������_{��
2����	c�f��eKU�c@�-5�o���¶c����P��U������ez�x��t�0��L��E�����D۳pT���j	�����7J+��5�ѭ`�dOn�X�5�; �-O�٥ٖNG���������F��?��������=c�P��L���	9m�������� 6��E�BJ�qY�w!%���"��+T<ק����z����xS}�����r�4{�-��]���{��#��T�B(�Ns$�Iԓk�Bqw�i
H���Y^*�m��I����}��@X�� �g�f��� �݈��30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�+ڜ4X{^�wLРr�A�}���Jdq��B�Ϥ!>m�gخ���T����r�2����,����.��km�EZ2�X�?C��>T�Gt�U�����Z_4�ӫ;�T���u!U�Gip�L��C��S��S��!
,/�0
Tf���3�^C�Q�$�Ť�^��!9]�f`ay�ȳkrMX�6Q.��� �1�F�j���xߖ��0�Q�:��澀��MN2�x�^/hĔZԙ^�F���[�J`�&�/�]F��M8^q�-�Q�H����2��:Y}�Ц�����л��8"�b��G��Z�*y�p�]����*b2yso�Ũn�U7w�-��h=*�a����<Wr�ۤ�f�{�����w�i�|N� �y��ZQu����]o)GK�Oz�::��S?SۻQԼb�a��#�fϢZ2+�jK,%��p>Ïi1���$��28Rc�"�	�+�*�ӻI��ZQ�X㷶G��F���O{"�>��-���t�<_⑽�6㈒6h�@5|����T��L��q<w��A�,�ʂ
���Y�J�+�������;�	'~��ܸ�����J`�le\^���"�ʚ�QٗS�.��O�XoT(�.Xq�042�¤�9BIdЁ6I��@8�Ӂ_6�q������C����K�s�L�H1��م�h9K�,/�6X����!��Kz��������B\��%�z�f�7)X*�{}x����6�I��f���DAc%�����[��P������ I���u�T��ē�3cr�%�Y�-�?��0j���Q�����[�ٹ�̚�Su�EK�h_���r�}��Bf_m�.�� �`?bu�~��*��W�:r$�s�f\IKs9mx8�ڗ�)�����a��v���t8U�XU�ľ�A�ҒR�J�����4��R-�Ա=��/�*��U����[Rb^�_Q7^zF�g<V�&G�-X�,9������t����.�g{�l�:N����lT�AG�ntk����9�S>�£~�ZB)/��YA��a��V�	$R������ �õ4�������9(�O�:K�٠S��m#�2,�.��476�&(9
Ma����	$������c����/.�<���/�CƎP0Ϣ�P��)�⬔�5�"�N�=3��eܨ(�����ϟfbԜ��!��``]��D�Yj����b����'UnMF�Ma�>6Ɩ�o�,�{����]${�Bv��p��}���76:�R�}�HcT�g2�@���-1���J��V�^�ܔ�D�]����[5v��Wh���k"��z� ��˥��]xm"�y�/���.��7��v��S���O��E�ӫ�����D(x�eڵ7���<�c'���Ƚ'��Ek��X�D������.�µo����,��)���|V�.�4�b���F6��\Ϟ�S惴0���m������߭�;r��p��=
�F������.N@��u
I�����@zR��3�XAŅ䗊AҌ��@�/�56G �Y6Ri
-����d�mc\�F��������Y? ��P�0�By���:aiL��Q���>��D�V�Ggp�2y�g��h��K�ʴ����S�zTm'Q1���To�N��7w^e`�S��#�S�J��d��%)�d@"2-��Lnp��`�C�3�[Qw�F�����[�-5��k2K�E�w�kC�'� ��$�T��� �.y�kns"wG5<S0�1f`�$Y�<��Ψ���茢[a2�����A���bn��UϘ��� �&K����62�\��) ��C��n�ASe�k�k,��A��Ȱ|�i�oȻR�@��5�_��8*����Q�"�Ȗ!U�r��Z,��$"ʎ�hp����Z:�g-��f@��o�)��x�/"�R��0�4n���|F�t���o%��t֤G� f ��I�p:
���|�p�!���s>��:���.�71f�Iq���n�hX�tR�#C�$����j�����|%%08��� ��#T˨��&u�#�4�m��H�>E�0��U��e�C�!4z���kG"�M����qτ�h΄���Y��Xw�+�{�����	�I�;�I�䅬�%�y��U�ܼn�)�lh��r���r��*���Ǩ}v��U	��>o�ٟ9������_�.����q{\��@f>k��#֯QP��Mo&�}�/o9����i$z�����y�(e�A��� ���g���Y*o]��s�F���'�e�*���7L�<69�M?�b������8W�N��ףE�?L5m�Z~?*uD����1�/��ex����L_*��K�i�%cj�G�,�zK��h��^��_�9j�wO�ř�f/��^��6\�c	^�@
� �x�Y��jLx��E����&��=%'�) 5��%ؿX�8�6�܈Z
�z;8��XuĒu}K��R��]w!�L�&(� Zb-����l$U~k�Tg��ͮ槡���P��j��80�8�r`%B��ٴf�>Y@F�O�%���]�o�y��$��4yS)N_ҹ�[/r\���~G��/ A[�?˗�hn�v	V[��A��q�> olz��5�6vL/h�b����q�Y���=nA�ؒw5e���b:+�L�_n��l=�}e'9r�Թ�sZ���<�=J6=�v��an񑠠�E��ڪϨ4�9���Ҕ��M���vᝅ��A�f�.G����:ku�����v�=[GWֈ�fg���е��qR�#ù �H�t�9PԢM͝8(M�.���#�w��
ab�H����*����9%�#��b��oB)vn�%�w�
����5*	9�1�Y<��V����7�6��w$/�|�p��᭜�>�Q�4�j-U��Q&)y�������p��<��?�o�Q<����#X���¡�+R �,zg����������K��0	-8mU���_7+��N�S�!}%!&<;`އ9F��r8�g�]-�?�4��)4�$��0�si����Z��#���ē�j2�� ��`��{����7�4Q8C/L��R���_��ɶ��G�1�gWp�4��:��zt�������ߴ~��]��lF&ԧ�Ca��9����T��ĳ
�+��н�`.�F�q�+ �Xy)�w
-٠���A�{���#"˗��UW�C�m�P��C�ܠ�ˡ�)��2�.���I�w^[�Y��m�L�2?n?�U�>O��GrRoȝ�a�o(�_r�j(����]T2�u_A�Gg�LS�(��ؑv�!o;�T���q[c���ƨ�C���ӕ!7�{f���FL.r��m�4����!���}��E(�!��TQ,IJ��˛���@�`�OM�w
�E��x#�v�ZRU�-�\g�����bk�C�sA�b��� �(|Ʀ���S�\0��bK��Ǻj�to�������I�ݛ���0!`�I�\�S�@£�EB�J��2�Z�a��N�s�-����w����\?���[f��ڗ�*c�3Xd}
gC�s��V�($RwGk�p3���c�c�ܵG'&t��`=n�S~��pA���r�!�|a�v���q3���=��$� ��h�Y�_e�*�ʖM{/s]��42O{6M�$A�EH�VjZ�i�i�)�b\�����3J$���*]Ҷ�(�<�~
g��<����Í63�>����B�c���̳_~F͚c�쐡\M�9�nت�y�D��YP-؏3Q��^��d��*\�ؠX����xj�'Xɭ��2����#�Fy�j�SwG	�v�Qf H jP2R$����Dj�-�'X�p03�d�� ���Ѳ��s@3Yuq�s���j�1/#(q����q���bG5'�Y�����+��5� d3Q�4Z$i�&���Z����g���@����
3rex��p}����D�T��N���@p1e{�K�C��1$�1���A{{����҈x[�����@��2�hw��}�Y�3���/Kk���,��
��,�q��B�9��4x��B��w�8b�a#Ι�슆r��e)j�N�������l��:��d�K]�5�:��p��N�}U3J��`�}u����1�I�A�Cæ ��w�Y�.��e}u�K ��&��q�ͧ�:����
��;��vu1�b:c�G&l�FUŦO9�U�E�zSg<�%��-a�\�-}��O��T��!�I���
�)�����3\Y���Y%�㰖�ǡ�� v}�)R��n�j��C�z)A�����{��q��
}ȹ���X@��qs����V�(�U����2Bݣ�^�<_ 5D?��&N)a��j���K,�C���ࢭ�����i��J˽8��j$9�ϴ�<|�7�`WĞS�Y$���&�Y�	=�^HD1����R�����i�	�V�k�5ָ������A��@�֜�c�,<�e�7k]& l�N���;w/0���OC��x�& �`-k6�����@��|�ZfE����Nx~���P�
��i'j&�O�ɳ,�E���
hQGŤ��b�qz�2�ҟ�7���䟐_�y�,���M6-L�$@,<q�ڇ����ﺇe�,��AѠ�k�x��TOʆ#`��v�>�lgB>���RDJ9=Ӗ���S�粠k�l���.c���>����n���W�XU+%\�R�F~$�^m��v����ir�Q�]��:Sn�����Y�jr�(�<a�~2](��)
Q�W:��z��M�L3�hߔ퐢������ɌF� �s��U �a3Q�"�Ԓ���9մ,&�u�C.����O��ga������3�M_�.Ҿ;@>o<*c_�?w��W �qh~sH�q��r�;���c����L?=wd5V���H��m��y�B�|9~���d��}Z�G!��,��#��������p�S&��F����ھS�n��g?���;�=���A��c�)M��oȊ�������y�O�	m�z
V
�/�7�6�G�@DWS�!f�����Y�<�p��V��;lzBhO�W���˰.GQ牄��=A(BXa��R��7}�R��
�|�5�,�B,���O&
�X���ʙ}���B7m�O{:�NK^W�M]��h
��'o�� �߻�,Pd��+�k��W�D�\�@u�j{��%��1�����d�x�	����Ń�oOr��c�@5�1]T�v=1j��^ �['5V�!QH�\�J�LDk�L�I&T�˳�\������]NOe�����&~��\?=⇄����	���r��vS��\�q���+�B�T��S]�1��@L��r�מ���v#�A�̫�L���0L�������P�|���9�Z�(�UnqO'^�W�=�#8&����s��� �8Zk�ǆ�#��s��]tM�%&�58�8Wg_���r�! !�s=�8��H�)�"��^�M^w��}k������O�q��������-�M�\�O5zi�$m�'�7��*�;ژ-�?�=������N�4�L^UC0'�d,��y!O���(�$����4]�����=[ͥ\��,���+��fF�N!ӟPR 9��E���Ć�x؊s�Dޠ��l��c��d���qNێ%H`m4E-u���d��a����h�j����!z�Y'��^�B�dj#_`��\��z����!Q熸IG��y��B�ꋧ?�T���� ��Zy�������_h�$�: '� iF��*�nܜ�ĕAk�F./p�{J����W��i=�����;�> �L�}C�D�Ck�K8��͞��x'�OP�s"�FyCP���[�u�0��T���"^��|P��Au�Oz�1s�AԭN�����o�Tz����8�������x77q�?��8�.���[��>Z��%}���:z���I�`� ��3'ϒ�j��3u�?��6[u	�7^s�	���F��Cp>���2
"	aƫh�h�`�^��sC~��p����V�2�cTaY�=���lG0�Y-�[���Aw녴�0�'�I�95��s9�JK�T�,\�շ��纅]CJ�Z�W��XV1��_���e)v;�fw��8$,�Ձ�l���٘_$+�d��[�{���W�
9�~6���l��7�aN0���>��'�9X�~by�̥�5"�"�OG�I�BP������Ϗ��0^� �Jx����#����+~e��	$J�����.��1 I�EpV3��Jd�ycz.ڨ[�|�������q���u����]H[Ez�2�x䚌�+h��Ԩ_������}]��9j���?X���^��b���Q�y8�~f�W"Ev �.zU��aС��s��	��ִ{K�%|��.fH8/�9@m6_{�o�"�=)V{4y� ��:��`���UOO���X��Ж��Fi�HXy�6��!<��@$Ur<��'3'F^&jޜ/���l��eJG�r��E�C�j�7<��]�}�/G��407:��CG�H��	��,����<A��\���T�T$�%b|��	3�\N�����n,Z�0�� 
�c�V��]U{/z��z���5�A�)�H�J9p�٢hum�5~B���fH�Db+����v���S�7(���J�� +i�OՂJ�m����.�}�;���LJ��y\�����ʤ�	�Ŏ�Ǘ��朖��Ō|(���qI]�2Zc��E�I�Y�6v��a��@�_C�q�@'�ٶCl���Z��K��L��D��0㟭����/`[NX�������K�K�Г�i�,\�A%��Jf��X�4}"���'I���X�4�Q �%����Dd�=���b}���O؀�겈�k����@��c�8��v�-����)=�m?�QiSf�����fZO�$C��α�V��\X}a��f���;ڮ�͘��a�k'I*G��g87�@�&fpa&K���x����X��yIa���o�8"�s�w���D�s�S���撅��L0RZ �
Kw��6���ZZuR�_�~�^2eg.������:Bf,���� t���7W�gC��l��͹|7K�y�'A���_�tX�jW	k0叠�����/�N�AC���?��[𒣫qQF}Wm.�S�'����B����(�:,�����e� �m�f8,�����6F�U(&I6M����O���O��c"����,1��O��������lP����O���B����3�`�ܕ���31������i! �1`j���j	o�O~�N�8nz�M.�e63���|���(��@�-{����o�E���˄��N6�ZW�;H�bg;1���.1|c�Ji����b�����]z�؞�����D}��<"=���GP��r�˲ʘ]%��"���/�Zn.���7�_v��J�ZM�O�Uo��3 �x�D�e��=7�)%<������ʪq_*}�#�*D������[]a�<���4��i�~KVC���	�Ab�
��s��ӱ:�jc���-A�M-�ijD��ݧ������AVpm�=w���o/ş��{�m��%Q�An�֚���R2�3��C�2=銎@	��x���d\�b� �&�R�p;���dv#��f��b��|�֟/f�&�'�V��0�3/y<��:��m��~SQg��>����j]Z��g}PyC����oK���X�S���T:kd�I�aھ�L`7���`���5MvS�jkػ%ѥ��dMJ�-5��n�]`��h�zr���QD��	��#@o-������2�����T�Ĉ��j�����V��\�k�̳d�5�3}	$O-,Y*nr��6�)͢��z�#������n����n3�ϥ��x�9&��i��cm2u���V�\���nA� Sr��'���ޅȝ�i9�e�@zr����E�s�:���o3ȃ:���uZYl����"}o�������ZS��g5^fͬ�o�l��E`�"�S��@�4���=J�|3�;���oRJt�ʂ�mE� ��`IG�O
%T|�>!@m��;���U�@+�7>�iIoӎ�9��5�f#p��$W,��T.���UK�:|�cy0%|ѭ�#��Ȩ�^�uZ4�q.����>��40�i�U\��B׈!��`:"kT�q�����]�
�q)�V�׆>�XDl��k���E��+�;0[�r���V���q܉��)!�4h�J�t�br��n�T�evA�U�OX>�p8�F�N�3�W��A���(�������t>�l)#�dOP�'os�%19�%^��NNG�݄�眆�\e��Ҧ$:�� ��(�b*��{��j򳢁�V�eȏ�*��>79��6Ƃ�?�w���_�#~W�7�ޣ�L"�kmN��?5�$D�ɱ�D,��<�L׳�77LLTE��:��R������}���^ߠ��&�jj���ψ�3+���<�C���+׍$ ��M�����}vxU�>E`f��:��Q'Az "��%eޡ�eѣ�}ғZwH�;E�u��W�F�p�ޞ��2�yVc(���Z�Kҿ�"lѠ^e���A���ZG��Ω���@���{]8=˂�Y�B���S��Y��vF��%Å�cdoo�Md��yƁAS�(�F��[\il\��/�k�E� ��?��h[ɨ	�Q�[%�?��8��@l�*�5���v�4h�>J�x�����Y�	ª���25�ѱ�e�/7���Ő�̉����'F:��f��s��{�%�nm=�|U^/:�@�kM�BV6�������r$d���{�/��y�d���لgE6qi+���HZ�ug	N��q5�1�@Ѓe�2uՕ�ᔶ�]�_��2�q���ӵ��F"�݁с��<�˼�A]o՝"^�P/~3.�67+2H�t�V�$�\O�{���ƛ�H�D߀�e���7��<�Ή��m��:���ҭ�rD����g�֥�����X�؋H��cb�T�V�J��ʌb����V��]�$�4n�ˑ������3��=���O���p���=AAx��=����8 ���R��� ���w�RАz3���|v���ȗ�,����~���& #�R��Ϸ���d�3�լ�?b͆���y�0��
E� ��0�?�y�Z�:8%�X��Qq�>��6Eր$�qg�Ʋy�7�?=K���bRVS���T���hP��k�]E.�7N˶`P[f?":S8��Eeޥ\4qdW�-E�nGRg`N}���)�Q�<���(�-�P-���Bm���;�����*�A牺�F�u3�%<hkE��.dn5�FCS�����Y��参�Ӳ��2j	�'b��x����T�3�`n�Wϯ�@���&"���V2�����H���cn��S|�bv�e��g.iCX�����@.G���O�˕�v���i�M���	A�Z��c�tqJ"G�n�O���xZ�ލg��f�сo�2�����"�`*���n4�Z�ǎ�|�������o�stt-D��7�) ���I�dm
�S"|W>�!Jf��Uk��K�
 �7H^�Ih���t�jb���~?#�e$�y��-5��-����SfW0�Vѷ�m#�?K�2��u��4�����P>�	0��nUf<D�!��E�*��k^�,�D���� �;������� \X�w䊲��\t�@�;�?��<]Z�a��U��x`)�5h��_��(rwd2�~j��^�v�)�U`/T>�A��P���}��6�Ճq�O�ËC���=�>�g�#��P���o�n���t�9�n��<���=^�N윐��e�ts��mꘜ�c�2K�*��~����}��~e�\*b8�7k96П�?�F�<'��}6W����ԗ�HL�q�mX�?�Dj;%�ϒ�F�b\T���<�LLo��+Qޜ�<��vL��p�����^i���jtwu�<����pT����MOƸZ_V�� N(r�������x��qE*�p�@��4���%n �R^%o!�����ZA��;OX��O���L`�:�%��kM���(��Z�����0�lpT�GX�l7�dJ-��0.<���8GC�i��B||��}Y�C&F�%M]�--�o�/��������S��-�P�_[�!0\T�<������ 8��?�sh%�	��6[o`4�]˸�u]�l��5�,v#��h��Ս#����Yn�t4�ｾ5��������������9�iLt´P)'P�K԰t�s1�N�� =�&"�)g�Wa�#��l��)������+�;�����k�v��	W��]��.��?"s:�>M�8��Z�:v�Ǻ[^��V�����l�"q���0�SHL��1AJԹ;�/���\���S �7,b��.�D�*R O���Qbq�~o��n��Jwv�~�'d*@��H�C<����������� w���|"�����<Q���A���|q�)��q�<���O�s�?���Q3�C��n�#i��Y_�+�p�,�� �8I��h�B�A\�8$-ٍ��+b͹����}\�,<R�<�b�FX�8z��]��hʫH)�Ѿ�+)os��\��ʫD�׀ �����w�_`Vw]�;�7��]+�+:]CTz�	��*�߄U��#c(1���p�ι1�tzK���h��T��~B�]�BF?�Y�
���x0����A�NU;
����jl��FÅp+/�yXp'sw��M�KL�A�2���y=�����Z��m�U�pР��	���?25���A���� ��ps�m�XT2V��?x;�>�~�G�Z�����B_��|;׫�q4T�ʘu���Gޚ6L�S�O�ب��!������T�5��F��-F�f���z%��1[!.��f�!����kr";R���o��p��P���ʙ�I��+?8�J�&�� ��_�M}���#�oRxM��	--<Қ.���g�Rb�5�C�F����p�o��5�:\L��	�0�wb����drtf%�����8�j�2ǯ�Ӵ��+.d@��_�<�.J����w(a-�/N5��-Ea&Zw���SW/�Ǟ[�,�.66cE"�d��?z9d����(�"G���p�bپc�s��eCl�~ֺt�z�=e��~�a�p�0�	S+��[a�M�hë��8=��|�k�G���X���}�͊]/�A�+��{��$��E��r�)��iFJ��yg���|7�
w/$z�I��|�V�ŕ���~A2$�Sײ��896
�Xì:5B�dR�N u�
�!~}�}c0,2���=��n�a�yQ�ˇ�7P�f/j]��ߣ�����>��WuN�U}jqN���j2�7�⏎�=�j��w��cv3aWݭ p�W2�|����Da6w���ӌ'�$�������݁�����5�Y\�
挑��1��&�j��Q�	��LGLC�Y�#Y���u+�����f�3�_�4��������������+�@I�[�S�3�.��i�ű�Dܾ���uN�16@'�'e[Һ�L1{/_�E{�E��n@�_�Fߵ=���ȟ�
ohΨX��9��J͸���KB"�ƀ:����>�#p�9��1x
�����
�n�?Z�:��錰e��7N�������c���!M������������N���3a�`�M��ޣ����I������ �i�sm���u�"��v܋�f�2�>��:t:?�a]��/�㲆�u(Ԉ::��Gݣ�F��bO���М�P�gS��m���+\֫~}��\O-kT�-������a)�yr��\�6��Z���ж3ʺ�m)I��nq����p^z�d�#�N�q�'�ٛ!$Ȱ��/yhŁ�L���/H��FU�B��pݚ���ޞ1�5۰d�����Uj��KC���������t��p�K����8�+�j[*��Ff|�F�7��U�g���o�&ٗ� [�	t�H[�Α���RԲ��w�~ispGV<��5-!�m��k���]� 5���d�?k�ZL����o��r-+��/�q|X����KZ=�ЦE��� \��%�Q�fd�X
��}X�:��}ZI�
 �˅��$��%З/����0�>��ʒ��G����c�u@��su�cR���(�-�����7� ���ᨽ�،͖M��R]���~�	��r�|\љ�a:;t�����r΋|�+�~nχy���_P:Gȇ�1.yL�e�PG~��W���Ї�X���4�/b��|�a�4<"�/˔��\9��&����YcOۄ�a^�ڦ-�%3>��jh;���<fx>�F�8�'�P ~M3��Hc,C��;�B��O�ߍ���L{� �fV�KHɛ�m�qW���9@����d������h���e��B�����"p݇�����H����S�5=�x�{B�������AsJ	�Am�ɬ;��(�RJɡ����Nm��nVƝ$�s�����N����|.�BԤ��dVZ�,;���h�S���?���Q#�����(~Ѹ��'����3}���'�8~�Q��B�y�VD
f��	�}`W"Bs�eO7��N�PPW��0��I
n��o2�܋��ۘd�z���.�W�zS\�-��&��a�>1�;��Bdz�	�ש�f��ի��a�L|��1�vB���6���~��-c�������������1��m�K��]
�A����z�&�W��.=���A��	ݬ�r�n�Sʢ��-sT��5۷��;.���}@��(r�>s��pӄ��#(�s�g$��Cr��M��5f�JS�P򐴙w�ZM����qN!�^xq�=�t^&m8���r��x��t�9kl>=�_�Zs��t��7&ъ[�A�8v�3W�j�I��!\�s���*���U��%M���߀g�Z�E��q�d3�|%v��1CMk���Rj6�z`/K'�A��f�w�T��?�H춢&���p4��`UP�'t"�,���yݳ���$��z��4N�Bn���\���Н��	.�ܣ���F��[�!R<o��}Q�z��45�s�8c�Sx��-W� c�� $k�J�`�eW-1A
�;ȵ�٥�.ii�&�(�zDO&�9fB���#�L��W�z2�ՇݣN�������IBp;��{VTL���<Z����'��}�e�2���� c�giU:*2R���cA�^�.�Y/�k���tW5��i���:�J=aK����X��D�\>g�9�K m &0�?P	�h�Yf	��9[]|��e��,�l��5�{v�UZh�ЍI������Y�i��op�Ɇ5�c��T>�P/����������"<�'~KԞ�ts�;�	ކ=�j����a�����Զ�T�r0��i�z��`��UTv���7La�KJ�.��w��0<:�8�m��EMv:]![�aE�s���J�$��k�qD��>H�^��d����0�� ޳�:�H~��e�Lb�W���*���.."�k�b)�ogs�n���wdr����*�;�v �<�U�ۑ�_��1��uw�+C|���ɆW���Q�ۀﰤ��Ef)>`'_����.���)}? �*Q!���N;z#}ˇ���+�&�,Z��}!S�<���0�k��T8���ٻ�+P�T�X�}�I�<�W�m�F��8�Z�]�ʙ٦)9����.�s�^��O�Y{=����/��e��`Uʒ�l@��^F�a�C�XZ�w�{X���rC����1j_pѶ�gz��R�A�Ց��~0I]���F��ǧ8UĹfsz�@=����
�W�pt��e_�F1Õ+]�FX^x�w�X���#A�����'1��e|1����mش��Ȭ��������2#����u��Z0۞�Cm���2տ?曀>�	G׵Ȣ�����_�x���ΫFJTW�Zu$A�G��-LX�ᙽd���Ф!��s��T	���6P��q}�� ��({��!v(f��/�k��rP�p��#Y���T�o��d����ف�Q�u�T�:�l��eI!Mq����]���wD-[0ǚbs�zUb��C��?� Y_��B�M�c�h�Q���[0�%�b�R����tT�pIS����`�J���ȴN����@�k�*c�J^%�@H�a[��N#[-�7A�\>w�K�AB��u�g[��*�\b c3��d��E�(��X$(	�uG��pX�WISQc�3�����It�[=S�L~�F�pf�ɕ7���=a��h�siP���e=�P�I%3-3
�h�/���;�/��O��{�;$f�sE;��e���i�gè�2��׭B��Š$������{�D���Aϧ~��w߁�{��w%6�����,B�d@�<&#̸J�~��c^�`��%9������(y���u�P2�E�$��A����B.�����C	��*j_p3ɲP2G���ѥ+l/j�NwlI�vaK��� �2��*�DO���+����Z�)ջx�a��}��WUn�ԮY��_�-Z��T�1�Q.ֶ���e�:LNGz0 YܶQ�j�+e��:{3���4_M��^p�>ٳ�s'�Y�@�[��/W3זh���s�3ͳD
H��o�N2�8@��{e@��ҨY31)c���v{�]�+,���#���D����h|�%�"q�x�̬�g1K�:��4�1�r�����?�9k`^x8B����~���\�(�h�!��,#e.��N6H��⫹�Q���f���	"����.�u_PNBŇ3��x`�BXcq֨�zIƢۛ�r{ �$�����B�u�%��$=Ũ�X��lЛ:bܙe�>-���1�u�4:���GK��F��O�o��J�t�@8g��8
����<\D>�}�c�OQ�T�љ��(��(U)����gӫ\~�QM��H�g��Զ�q,��)7�NnU!�hz����$� 붕�z�O�Ȟ����i�|�z��?È-�#U:]�s݈������5	�,���f��ja��Kqr�ݳ7��2����������"�8��Gj��m��&|��������I��������'	�N�H��g��>R�Q	���^i�r6V*��5�f�}hA�v���|�!�c�e4�*�6k�<�l�1[Y���/�0�E�O���x�=���k����ϊ��֪|�{E��Y� x��h�Uq
%bi,����h�q~�E���
�u����N@1G �7�1�DH�7�O䄐��u�,�L8M�?J~��$E�lqErϰY�3�ʠ{��,�o&�e��{wK�Y;0�������Q��>�^�wQ�J�TG���X2����k �;��m~�"���}ց3��Ӽ.�XZc*%�<�iQ�C�T�F��2����r.�<�bGL:�Y����>))r�Fa��~�W��"}�V~�:0�?�:#0L��뙢Ɣq�G���W�g�K�[�3��j�a��"ĺ��>9��&=�H/�>xO�k�a�_��v��3��a��;�P�</�E�/)�0�Q �.P���H���7��;N����ԍ� :L���I��VN�&H2�.m~��ڧ��9	G��kNg��xY,�ڱj-�H��ˤ3�d~p�QS������
S�����j�!j����A\1C�J1�Հۊq�S��}��>�Ǝn _m��V�]'�|p�,���9L�F����B���k�u��VC'�;�l�h4)r�'$-�SϧQ���Oc(G*������}���pW������ڭ�B��:�V
O@#���}� 4B�n�O�l NՃWU����p
W��o; �N���Id!k\�0,�WZ)c\������j��1�KT�d�T|	SN��?��t��Jʁ�p�1B�\v�]�V5F�|��Hj�,��ƌr�����1���w�K�͹����GԐ�U]�_��21壱-&C���=�Ǜ����	��r��%S� ��V��6Z�gǗ�Ĉ��ǭ@Qor�x}���$��
�#q6���*����I������?�3f*P� 홠FcZ�w��z�q�mc^!O�=��&V$���{��޽� k�����sA�=tR�&�O��8�J!W�r�����!�)Ls���������t�B�M����F���}Y�㔁�Wzq�";�e�u��1M���!�=����_�'H���/I��=��?�
��ߐҋC��4���U�*�'�s,���y��1��I���"�P�4����ː]Ƣ�եa�����������F`�S��}�R�
�۪�t����s�p��|�K�v�7艊��8���Đ`r��-����l��+x�w �菆q���z퍷� B�F�#�v
�Az{g�F}��}��ip�~�BY����)�Tu���c~�� �U�H�&	�������� l�qi+�*{������A0W.�c������ �W>��i"�a�r��;$ji��C�sD�����m���	�� 'qߐP������C��N����q���@����=���W�åⳁV����o����8�x��T�wk���(�[����^3%0���M.��UcIk��:���Ƭ���j������M�u|ց^F̒����ѥg�c�{�!�"�dP�{"3��Ο^b �C��ap5�X�I�븶�1YpDt��I(0-�)�.%+�t��G�������T��&C0J^����nN~f��"�G��neJ�W�EV��o_�<A��.q��w��
$� 1���lH���S_71�d&�r�N����^�9$Vw��wjlf��7Jy�t�h�zz���z'-O�9�6~U�aw[��7@5[���m ��l&�b-��#�u ޘ��=6�
��<Ze�h$}0��\fz.ݎ� ���E#r����uDN�z=g[:W��i��à�
]�����R�Hw�zy��߫$]����+[�9���H�X�cǐ�	̬�8��XKi}�� b4 �-,Ry��f�XE�=�.M!��էz���淪Vs(����{^�"|��.97�b{�@ �_n���u�)	B7{G�J :����ͼ��\�U�!.�����}��t(�,�yj���p�s�XU����'r��&</������T�=G����؉l�]�s<K�]��b/Z[�4�#h�e�2�{_ 	/u���w9<e���	�g����d������[;	�P�N���/�sZ�Xa���b������{bUƨ(W�(���|�Ǒ�u��Ȭ�h袕5Q&��Ċ�׆������
vl�/�J^�� ��JX�J+DJ���	��=�5�I1���.,�N1���J�/�����\��m��$��
���A㚗��"�	rs�٧(�q�*2M�x���I���6�����,P_v^q[�J��y�C�ٖ���KκL������Қ��0/Sa�X����aM*K�p��兝<�\6�%=5�f�9ZXj��}�sb�#wI
ϲ+q����\%0�&�7��������;l�����[����t���c��:$�-^�<�#�O�Q<r��,�!��y)�a$P�������}Ԅ�f�EL�nV��`��d���*�F��zLʴ�8fC��K��xx�c��kJ��na6h8��p8�������"��Q�F̓�9�8�t�JRm�f�}g�o}��4�T��R� *_H[4^��5gA־�P����mʠ,y>����t�H�����gVUl&]��O(z��5A��R�4t�1�Ĵn��Κ�/��sA����&q.!\�VVd��ʕ��&�˳�<������(3���zf�����hmc�C,7�1�W�;69�(yT0M�@3�&{ad��"g�cU�(�*i�|ʆ�o@&��"d�⢾P\��"W2�u�u����3�S>�������������9w!ӛ$`��-��d�j�Q�ܢ�zen���M�Ƭ6���>����O�3`9{�+�"���I�P��6zc#�/�H�NTgr�S���1/�҃.e[h�՞����6{]9����ǐ("�=�&"PrŁ����E�����3]���"�;�/��.SR7�@j�]���-�=O���ft���vDh�,eSl�7�m�<�l��l���٦�?X��hD
u��Us��n#��f���b�����V6���\��b_�L놐��F���=>܃�b\����\��1��S���߮�p���=J
���'z�2M�nPG�G�\J���j�逜TR�R�3�
����݊���˚�Gj�uP� ��R���֦�d	��}��WW��/�ßB�b����);�0�t�y�4:�+���QP�>�y�.��-rvg�My�!���wK5��MS�T�T�I�q���!T�z�7���`��-���S*\�.�٥e��d�i-��an���`�?��%��Q�w��ܔ�V�-C�������
����gq�*�u���`/'t�n3�k�u�Q`5|�r���TY����[C�ㄢ��))���N�������an�p��Ȋ�[&��Kq2(o �iz��$�n,LS�ʀ��џ�P|����i��u��vY@��[�x�B��Ql�b����k�C�Zl�[�]�M"P4�7k�0��ZF|1gm+'f�m�o�C��w"�ǅ��"74D���0��|�Q�8�eoe=MtG��@P\ �,\I��
��|�z�!�3E�ر�z�b�Y�7q��I�]���p�벣���#��b$�.��'л%���8��g0x���`��#�4h�$gu��4�_��B��>�'<0F��U�v�U�!t��3�zk�T���\��PK������(יg�X��h��%��/:����;#L ����e,��0�����)�֎h߉߱�r�Ɍ�}Q�{yvToUI!�>�p?�y�5�����_σ�y���&�jΌ��>��P#�ZP6K}of���oy9E{�����W?����_e(�5����%��y�*��U��%��B�Gًe[y2*�z7�a�6yg?�|%�%u�����W��?Ω��jYLu�\mm?H�ZDSj�����o(�� �*�L�4|�%��e�%��~[��u���L?^҅��yf,j
/�t���Q������v븣׀L� �顙���tx�~�E3~sY�}_R�� u��%Ҕ�x;���~ZJ�8;xIQ͘勒�?\��\����k��#�(�'Z��Q��:ld�,X�:���`�A��ْ�s����z8pfP��Z3B����A�Y��4F�i�%6{�6�o�kg�A^��t��Si�����[o_	\=�=i�F�� ��&?Zwh��8	^TY[8W��F���~*�l�N�5CLgv�1Yh4ڪ��}���\�YWǕ�}�$�E�5F_����km[2�>���R�Z½�'yd����s�-$�=�H���PKra�ہ��%3�/n�k7DP��$Q���;�T�.v!���2)]��-.��޻�/�:F��H�U�C�v�q9[�	`��`'�O���U�q�q���vH5�1:�2��?�xb��n��cS%���b[ߑ�-�C*!��)lK�ch�b��io�3jn6x&w?����H*Ic��q)�<�}9�L߄#���v#�wd	�|����!���jQ/��o���f)��::X�����|U�?�a�Q|��	�'#�Lޢ�+�Z�,�	�����7:��ECp�!8�_1�6�e++pG���-}eK�<{��BuF��%8�]mO��tc)t��4��s�^����fZ�	Om֪��@�`?%��DD4��)��t� CoΧ��w�qx�M#����1R�pgR�zouz��+�\�Α�1�~��]�mqFHPu�3�'���I��Ȁ��`
/�דK����PcF���+X�X�#iwJo��~GAK�?���ab-��  ���Ԛm3�ˮ�NE���i�e2���*}���H�ۙ��m���2�U?`�>�4�G�����_��R�_�jZ�p�Trh9u��nG��tL���X)i��(!Hi_�.�TT$L��-��L
��O(���X��ű!w�f^d��@r˻��t[���&z��|��w2�V�GߔڰlS������NĀ��FM����ո����x���-������PÆb�S5C�%��[\��D�hk��A���L0�y�b�.���\t�"�MS��������p{洉F�>=@�Z����J��[d�a�L1N�!-.��/�w�0�����0��[�u��L�c�d�,5�;���(dLMGO�lps}�Ĉ�c_-�N�ȵ�ўt���=�ٟ~Xl�p�n<����a8�a���\ҫ�:&=9d�2@�R��$����j���w�/�χ�t�G{vO�$�d�E�Qp�����]iO0ը���2	�s�$���j/z�C��|{�~J*�|�t�1�26s!��5v�BT��b���G~��RcY���֨�y�9��@y(�\�P�Pm�qs.o�<�ʥ��j^g��~��[Kj:}���2���u��sTj^A�w��	v�ر�� Y�.2��3����D��+�X���������S���`E���r!YP�%>6�u�1oue�I��:T����Gu��Y7?a�%��+5x�@��3���4�F"�����9a���H	�@�Q����#3�̸��T��X�DG��MuN�g'@��?e��3҃�s1drg�%�+{��D5���:�>��ހ����Ch��Ś�ҩ�s�ܬO�3K���Ov�1���l�H�eX9-+x3�����xG����o��]����ei��N�ٯ����)xH�u��k���֛zn�����N�gX3��]`,���Ш)<�IA�]@ �jD��=�u.]��(������:=�_�J��٥��۽ruq��:�[�Gf��F��2Oy�[Ѕ�Y$Ig|fe��m�\_wn}-�EO�<)T�8I��w6�#={)���"`�\��Yȫ��#K	����<+���|)�]Fn�l
��.zi�Y�fj7���0�ޛJ������瘂`��F���.�,5�h"�UՕ��$&����BA����5�Q�f�����j���Kl��E���C���(�����e	8�s>jdc8��,=|���=�ޝ�噶/�� R��{�	}�H���Hz,R= �� �si��V��5H�!��^��zZ��4�c���⥥k��Nl-�&�0{�:07�UO���x(1��kv�)�F�S���|�̟E	�o�Qjx��ߝ���
 �Oig��ҏ?$�l��E�q
���/����rj���/^7݈���s�B�b,Ή�Mv �Y�!$��Nq���T5=�%���',ؗ������V���1{�c���3���!>O�_˒dJR���[�ԓ3��'k���(Z����{���Rfӗ\X�o�%����p������V���Mz�!�r	iQѝ^�:�XV��)��:�r��M|k�~r�t������:�)a�5�~LE��Tj0�-����2Ͷ��Јٳi���asK�"��fP9�U&���g��~7Oߞ/a��N�1�%3���n�;��H<jd��)�+� ��@H�{=�U�;)���SE4�'�L�[�ŧV	רHM/�m�u�ڂ[B9D���M���=�l���c=��F���^��p�Ţ&��r���2S����1��j�{���!�A���E[<�0Ꝋ,�c�֩ ��A�I��m�\�VJH�weTɇ��Y��a�'������ۤ�_V�Sk;�,�h��Y����n�|Q'\�*X6(����"1���)S}���+�h�����U>SBl/��Z�
�B����}�-Bw/�O�D�N���W0��K�
�%Yo6Av`���.d<.h��RvW5l\�b詪��eo�1^��+Jd��	ο���Qկ���P�'Z1���vF�q�r��pB#�fg�E�a;,���Ќ���d�f���>� o{]�y�����z&������="�ń,	��2r=TgS�8Z��̪�\^��!�?&j�q�@��/r-h[�����M�#,���o��G�Ŀ^���93����P��M����ZQ�̕VqR�^���=��&��u���;�"���x\�k���c$sׇt��&U���A8�EW��\����!`�s}ָ�.��i��Q�MT�����U��nA�^�g��"q�A�� �ֻ�_�M��J���s&d�j'#Ҙ�js���WU?����:�ԋ�P�4�eUT� '��f, 3>ya�ʸ���	e�]4�uh�F�o�}u&���j�lS����QBFф���R@K�ۅٝ�#ga��¹s�v��v��1&d���$ĩ�ο`��-�G��=��]�2���S��z�3�=��B4ϥ#�h��ݕz6�I�a�M���D�8�FYB�����XT��0�@u���C�����6<�do� g0Fi�c�*617��HA�[.o
��,Z�W�uW9�;i}Pٮ-��;?�9����C_]�D*f����S�Q�%��',�P��!�XjC���țI�p�3T��Oɰ^P�P��Gu'b9�q�+AP��x[�����}\� ���x�<���Q�Ձcxwܪ��xۼ��[�����%�%��zT���@I؂͈G���s!@�ЬL���ڽ��P?uI?�^�N]���R9+������"Is>��㬠�K^Ͽ�C��p�'�����^FY�����0�;����~���Ѕ�?��g�T�yݳ�{J�h��ZN��?>�/��GWJ;��W k�Vq�M_׳�ो�{w�w��:$KfY��l	�R���_d��d����2���9��,��o�lS�ĉB���Y�G��~ }':�)9���~�{TN��u�bbi���Ƃ�N��g����p�X ��B�˥c���ȍ�e7m�$����	 &.*~� ��mE�h���zn�T[ ���D
ײ寰��Ҍ�U��H�HD=�z�\.߸V�0T+�����/��C-ǽ7�y� B�XXXv���bU��_yx�Sf�q�E��5.�����SD�MG���;s�ts��W{�1+|ݿ�.�2�o�@���_��'�b �)�i�{t� ߉�B拌�~U�	%�\�Έͭ�h#Jy7Y�a�eÀ�"U�6� j�'_�Z&��*/*�V�R�<��Ge<�+���p�<8�]"��/��4p���-%���@	�s.�?L<RK��Δ�d���k�e����u�	s�TNח����Z���$��䣼|�9�?{o,1����u�.�i�ޑ������h��:5��Z��X.����������@h��h�w�F�ͥ�JŅ�+Q��|/��k�6ˎn>��{2��ލJ0u���\K�K��2��Sf��/9���������()��q�W`2��s���I1,�6�������f�_��&q{$�9�C�����K.fkLڈ��<��߸8�/�qX��j��P�K��G���<�� �\C
}%�x�f�XW�5}E���Pc�Iԡ���Q���y%�{��TC�}t��Ok�<j���!��]n�s2ĀGc���'Am-���i���,Q�=��9��٦�[�d��
�5�<�G��}��f.u�{L#�S�����q�*�{ǳ�����7f��[K���x%�G�:����a���H�y8b�"��7���>"Γsr�&]��_pR�eB�J�ܼx�A������R��-_5��^G��gn3���H�8�z�,&jP�Q��t��w�dg��-l��׹������CA4���N�t����)�I�������2/�@�A������&��j�����Γy��	���Q��DVq( Er�F�~W�`�?mА�,D����6���(f�M.]M�S)�1(��T5cbC���&��\��\��[|d�.�P�L��aM���;'�3�0��k#�sC��)�ԩ��!@å`��ө1*jI�u܏]��M�n�%�Mn��6sЗ�٩h�&���{�?��T�꯬�
K6���Ѿ�HP��g�}���[Z1�5��[d��L����,]����:�����N�"}Ny����i����]eN"�/�d�.��(7!��*�a�w�O�����톛Fz�DU��e�p7�<�᷉3Bz�
]8�$�cgD�8u��֛wq�|?�NU��\G�S^V�(!�I_b����T���Mb�`�����ϩ,=�踙�H����p��&=�6������H���$�4p����u��M��RF�G3�C�r7ߊ΂���U��6k��7� و�RԷ��Od�]�責D,�ͼ��o�a�f+�񖾝0�e�y|G:�߬Έ�Q���>�M�Lf�g���y�����K	$Iʘy�S��(Tz�K޳�롌�;G�7`Ɖ�zi}U�����2!�4�,s�,�>�Ɠ0�8U��2�?�U!�@���zfk1+>�w/�zt�.*��nD�׃��X�e��%������s��;M�t�/�RU�+�&Ʉ)^�h�tܱ�+Ar
o�q_{����v>'�Us�u>x�#���SF��&	�d&�[���؝��Ta>a�#���P �o������9�G��#䷓���Мcbey�A����Xg���J*��i�$���pb���eE�*�f67�k�6#�l?����O_<�`��W�)d)����YLߵ�m��u?2[D}޶���X�9�����T1�L	���5���O���|�$9���6��^��.����j����{������� I踍��ת� A5�C: ���Rx�E����]��g9�DÄ ߢH%�[U�b���Z��u;"�2͂����˟-#�G]H�v,*(.xZ�����qlN-j��%��A�շ���,I�C#g��8ɽ��MB����Y*{�F�=%`�S���o�ع�+` ƞ�$S�<�ң�`[YFL\gn�l����\� k!�?5#Qh�K	�["�7�p� ��=ld�5-�v��Vh��R�nC����Y�����f���E50?+�9�����ܾu���|0��'�5'#����CJsĔ�S�=4"$���z7HaM���4�|��9\�Z������@}�~-�v����ѿ鐄�.�s��2#:����2o.�m�v?w�[1����h�/T��_ �q<iw���H_a���{Ԍ�g�b�=ޘ����ǻ��-bE��W��*�D��2M�Mb��o�q�n���w)&f�:H3*��Ǐ��<�c��v�����ͥ 9�wNԙ| ��ɋE*k��Q_�Ԝ�o��)c�$,�����L�?�FOQf�c�3<�#�[���N+|� ,�E ނyT����u	#��8����R+۰��6}���<%�@P'F�8m�z]���^V�)��璞�sSac���>�S�sI��TL0�*�`i���cC��6��^-uC������|}��7���6N'1o;�p�}4�d[�z�$���7ޑ���~�h]\8F����b��)��%��Ag�
�#��5�a��ȢF6Y'+�
X��,wt�6�>��A�%G��[W�/;�jGg�-	�mU]��U�|�F�/2�7��T	��!Zo�C�bm���2钡?k�>9�RG������.O_\N-D@��+�T���uIa�G�L��J���b�{{2!2X�X�bT����[���6�*�yR���3�"�!a�f����*3ru]�^2�� ۾�Y�œ��t�@��߾�'�1�y����o���iMv�h�(�բc.�4�G�-��6��Z��z�rb!�C����E,����x즍g�}�0̌b��QǤ�t�<�.�¼+P�݅���Zz���"����@�d��o @JC�L��j	a� /N�V�-Xz�9�w�����t�Zb�[��ځ*Oc��
d�g�0v���4(ND�Gy�p��np�cI���x�T��t���=��~���p�ҝ�\�PK_(a��x�ët�H=#������_R���jl��!�@�q/]���^��{���$�\�E2Wp����ui�M�L�o�)A���n$mTo�?R�	H`���~����&l��h�6��ß�B�*���O�.N~�h?c�$�ˊ������T�yҺ"�:��P�pOݩ������(�J�V���'j$���^12LG3����p�aj���w�}�v��G� ��w2�ݕ���ID�qO�x�����N�=P ��"�\y?]y�Y:�	h�K����1���
��d2��?�qG��Y!e��Of�+�V���G3{4Į��c����'���J�>v�@<d��H�3��X�%�k�8��D�kr��N__@�vee9F�m��1����{e�.9����ߨ`��*J!��� h��?�'�d���9��K�"���8�^�V�L�6��9p�x��u�Ǧ���%����F���>�e��NN;���#F��6r��p�GFU�d5Ԝ�>cNG��34�`$�H{d��
�I��mn� $�|��լ�8u|�	\��YTt͑<�:'���tn�Cc��(ru[��:�1G�XF?G�OcUЯ^mëDg&��O�賗*x\ɣS}�y�O�+T�i���O�ͻ�)�[l�L1 \�1rod����1�>��F�`x)|�[n�����z����a~�������Q������g�[��������|���U?El��j���l��	5�5.3E�P���}_jf]%Kg����1�=b�gp�ç�tƑ8���jΦ\Ϟ��|Է�ʆ��H���C���٫���'	�,�H.��2�#Rg-��jQni��0V�z5@���{��H��ԯ�̢c=s��O��k��2lW�^/ %x0!��O�۝x�w/��&k`+�p?���S|��E��>�wx(���:��
�i�����tm�q$E�
�ȗo	W����E��$�I/�7�u���L�l�%,8.�M R!Cw$�QqJ�9��+���ܺ�p,B�ъ+��@ý�����B�`4���7�>y����6J����VXԽ�k��zk�)�Έ۷w��9~�X��Ӂd�X�Q�%�4�0�@��Q'���F��z�r������,:�I���-��.r�[��&~\�眴��P:5原��cL/+��~e��;%�lՇ𡌰P����?0a]�"�锉�H9��R&�x�q�ͲO��a��ۦ[�L3,��f�;jO`<��r�4C��� ��ٯHQ:��\�;���}c����L) ��+�V3��H���m���l�.9nHy�p|x�gg�q��ږ���͏���]��HBpI�͢�h���{��S(��fN�)x^�e�X�&�oAa�1�����.ЊVN��@�ӡc�=�3��m��V�*��!�)�q������`�Ni��Ii��֚VH)!;V�>hy�ڇ����K�Q�#��(�p���8����}���U�s�&����BV6ۡ�շ
T��뷓�}΁�B�-O%S�N5��W9~�G�M
\Y0o��3JDv��d��U8W�:\[�����1H�'�0( dh�P	x�]������3��O�d*�1��.vpF�:��j��Q�㖾�̞�F�p�vRO�u��Rt��	���J�]�ԩjHZ��{y&�U��=�'�G�	�r�ySx�������뤶�=��[!�@��br�W�׈�F����#Vs��UT���ܿH��cgZ8zmP�����o�Z{�1��o�q��\^撼=��&[m3��u���ޢpkZ::�Z�s¸t�_�&��0��B8�]eW�7�:!
3�sg��X�L�Ӧ���U�M>2�����U+���yzq���j���nMٺQs�$�u�'�㨔Y_�Bv?��.�$΋(<4u�aU�2�'�	�,*��y�.�����5�U4�;����g�)���َ֒��J�FE���I��R�N�o���M딎"�]sw����˿[�������?~۸�q`�$�-�j�j~=�r��\:�r���z�n�gZB�ls#I]鵆}@z`�H�� �����.F��hVB^�N�)�&T����j�u�P��z����R�`���Π! ��ip�*`⎜~��AU�c.Y#��b���<W���ig�L�W��;�)��63CI�;DT&���gl۷��a�'VWrPVh���CzGN�œ��2�T�bD9ۦ^?��PD�	u�#B�[�LA>$[�Aҕ�YwX�ْ�*k����y.����x�w���"�)��g#[4ޢ%g��d��)FIBpш�Lu�]�����fP��)����%^us��^���&.�<s�7�xYR"�\��!U�ʰ^9AcCh��p̘���˸�Y��k��o0$���-l�+�g��2Ƒ&|��o,�]ɲJuҩ�^�UU���\��1o�Je��Wj%V��_��?��%>�V.w���$5���?��ls1��ü�_N�Td��%=��A�`9��M��
l�0�n����yb�q'���'�m�9���~�.�.���ULD��*������R ������� 5�Q����M�ۘ�OMe�t�������t`� �U���G�dcl�6��1���I=5��]�3n�[`0��y)��:;u(���bQ4h�>� ��̠gʩ�y0ZC�B��K��L�%\S*�TGʃK�(�02�l>7Qށ`�ΓS[���A1�?�d���-"w�nJ�
`�8���,�LN�QQ����ۛp�W-�u�E&�_��ŕ��t���i��n,I����SbkH�"��L5�_�vɊ:U�Y�"-�(RG�v��5�g,�h����W���'�n�D(��99�e�&%9�%�2B�u�ë��n��S�����a�j��ӹi����a�@��a˳g̒ԕ'Z*���}Ȱ�h�̥Zƅ:��"*��Q�4����Z���gG�f�I�o"��RdV"�eN�|4�$I�ʌ�|`L+�R5�o�Vot��R�(j ��$I4!�
��|��'!������j~7�%TIN�wl��!��.�#�.0$dg>��6�?�蒶�V]L0R.��zU|#�{2��Vzu�S�4��k���>{0 r	U)0¯��!I����k����z���4�Ϟ��������"XQޱ���Io5��~�;�/O�M^}�x�Tܖ��)�
�h�8�a~�rz����k�!'�v�10U�;�>��	��N� ;�97���D#˳�fS��>�70#0�/P�Q�o X&�I~�9_���_��T���1!1���e��������Ve���*	9ቔ.~�`'�apge��*eǗ7f�V6���?5�}��w8���rW�����*HLO�#m{�?�U�D�f���jЉ�r�t���q3Ly!��i޿�e�!u���?��!��~^l9T�S��j7I�_�@�@B`�x������ed��f �c��6��@�xbilE��-��{��S] OA3%2ȓ�����c�Z$�i;�������Oᥟ�1(��9���(��<Z|[�
(Fl�O��q�n�j�'+˧;\��K����D8��W��'B�$����Y�7nFAQ�%�M�.o�L���b���SC���ش[� &\�v�����`A� ۓ?��h�~�	x��[�����a+�X�]l�#�5���v&��h���O�rlY�p�W�W�2�U5��3��"�E�(L;��ϐ��.'�-��S�s4�,�q�=��EZ{���a�#���h�鉮b��������d��2+p��e�v�I.�L��� '(.!d%���:`�â����Z~v�-u[�@�({A������n�q��	�S�iH�y�������6��n��=����ʬb�P��;*��iC������bt+o\�.nP�|w�����@�*#���ή<Y�N��e���H ���1w��|�#L������Qw1<D�ʄ��M)�����|]��V3�?��Q��ꖣ�=#r���J�+�C,T�����?�Q+2��=
k8�Ԣ�P�+���-Q}?�"<��xrEF[�8�`�]����0�)m�'�   ^   Ĵ���	��Z �vi��:'��(3��H��R�
O�ظ2a$?�K&����4`��̏;Y�����,�P���#j��6��¦�޴J�������'��Ɲ����dL�KOZ��P*~�n��ѥ[�$K8O����7;�b�O�I� [�8IH����5�D5��I�=^�;�M�LyR��	�Ay���0��	D�+�t�т�/���`옅a��W�o*X��p$�j���Ċ�<j���^}b��"e��2d+!�ĕ(ǂ�1mȮ&�"��xrd0hK�yZD��tf@8=���2�'�9c��9E�8tp��с\
��O��"�(O���N>��&�8� t�d]��P�D��<��=��"<1�AD-0l��u�$FgN�i���j]�`���4L��I�V� ��P�W�\%��Ɓ"hi��'QjEEx�/�R��� ������=&�ć��1m�%��(�t��3%h�A���4��b��Ƞ@O�U��%5�	�bj������D��R$kx���ʲN��a�j�<i��5C-�㟰l�]���#�>�F�8wA�p>�t���	�n��,�|T�$XG��/$�4���'���DxrKc�I4/�t²*I?��\Q��*2r�ɩU���9E�Ʉ ��Y��"P��˦&B)nN2�Ę%n.���NS��3�a(�]�Jis0�.а���	n���E�L!^�l�+#Q���&o�0�H�Od�����?��'��D���L�(=f����t�8�g0��,zJ>yw�\���T�<��퇱 B��D� &@ܼ��%K�7�P��'�ղ@ ��G�!�$k� �  �                                                                                                                                                                                                                                                                                                                                                                                                                                      C  4  �  ?  �"  �(  *   Ĵ���	����Z�/C�'ll\�0�|r�'a�	�Dط8��0b�
�<�}#�'�t4��B�h�d�w,�:?������i"x�	�-��K����1Bʚ�HH�� Ҕz�J�[�.�0�|)`��u�(��dů,�HP9Q��#,��5˃ݕF4�,��	�a�l"�i_�6��	�aι ��0xЅ�)8���ڛZp2�"n�}����D�
�ZZ�Q�W��".ٲ�0V��	DWC[*~��?ѧ�ϔ&��g�WK��ؑ7�Lw؟��G�i��)p�ىH'N�1�Kò
�qK����B��B��};�6	Veg8D������O^��Eό�	0
)9O~���<���H"��^ӔA���QN�<	��A�<�>��t�)��"V˟F}�a݄cx0�J5�%��S�*h"`�5jO�2��	�uD	�w7B�bajE[G�Ď@�����L�8	�OLc���*m�]��ɤ!\��*ыUu��y�N�?O�:���K�	�B���гJ��4��~�0��Ǆ�B�	Qa��p�I�0��рg�
�"?	씛b����#�8'���ҫ̸X<�9o��yB�J�x��c��e�,���ܣ���H_�-�{���2�|M���T�x7��Za��1P!�$�3#���7��$��I ���%J�'�\\�f�Ix�p�Qǘ�$϶�@�O�ک�ҧ9�O�5ᄫ�1�����Ƅ�m�LS �ڵ&#Ш�ȓC@���VƇ�78JUQ�O�A��D~2%W�O϶�@o��*��ң���B�'ArA��^� yJWj�$D�^���'rf<r��O�Z�iw�C�@m���'�x�+�%S�t�G$�N�2�'��h��f&��ݥY�paS(2D�xI$k�X���yA �0j�lK�)5D�T$�K�m��0��28�딀���y��� �X�3sl޻b��D5�y��z�S��.n��isjO �y��B�m[rCU���\�KΟ�y�ɘ�����Џ�p�����Py�'��.��怛�)c�"�]�<1������q��I�:���QY�<�0���(�~ 8b[7e�m��,�X�<���vR:DY���fɖI�P��x�<Q���1��i�edH@�,]J�<10C�$b�89S �n�B���%
%D�ܹ�l*5d�x�w��l�pe��>D��#p�����- v����0D��k�U��T�����|mc��?D�0Ӧ'�9�
����B��(>D�|�$@ثg��@�E�*l ɛ&B)D�r1MF�s�ᴌ³ �<#%�6D�t�I�%&ԉ�gՖ��$��M4D��1S#� 7)���';��ՃVa0D�faR(:�4^�L�����B�	�2���@L"_��`��ڥ[��B� �|��	,p��PEÙ=�B�	4)�֩Z��8X��i#H�9��B�	h�OV?"x* ɐf�`ʢC䉛	�89�bC��00�@A)vB�*O�,i�,G��ԳQÀ�DJB�I[����g�4Y��C�K��! 2B� /��䉷L�57���sD�$L�B�ʢl�s� I�Ti �۫*FC�I;@��L���2?䜀 C��4�*C�	�[�:*�ȏ7+�xe�! �\�C�I�`@��iɄ$�T��s��%�0C�	�p>\&��%k�,��q,K�O�C䉋
̙iUg��t���j���C�	(>�ꭙ��U�u��QJ���,�C�I[�jh���:��	�V(�'j<8B�)� �DHG9&P�� �� =��"O��SQ�����c �	�"OB�c�gG�[�~h
 �Dh8�#"O`�A�L6��gfl��+w"O�9�ΐ}r�/��|#�n_2Vu!��L%~�.A�UHU�^Q�"��+kT!�d@���Ekg�B��Hrb�^�DR!�d�*�~����H��$Rc%�0(!�ā-[�d]Z0���9zAq���(L<!�N���@���%%D���`�P!!��8�@	�Ī�n�Ij��{2!�D_ +���A��4k>Kq"ؐ&!�D��y0P��M1eH,����N�p�!��2kr��z���dA�����:�!��/wSx��M�Z����5��	Q8!���}�p��#)_]�T�P�RM+!�٘fi~��.�.���i��V
KC!��b�
�Y ��B�nX3$��$.�!�ėua��0��#���*��"m!�D�5��X;7�1:�12��(?�!��`tȸ�v אN%�T
1�e�!�d 2����HڟY�e�'l�3~P!�$�!-�ԨhV���i఻�`ɿ"�!�Dr0};r�۷V"4[ �Y�E!��U�:�J�# �UAD�2�!�A6���&�.aը��k���!��NP8X!��[rĘ��F���!򤁃fr��ڇ�N#/O�|�Hާs2!��T�,��nO��cT��9V@!��,@n�5��훌#�֠8�M}�!�Ę�+D=��	Y�Q��Ղ�JՓ.+!�N�A4JA���P�W�b1�ႋ?.�!��9Q숈������L�D�!�DC�p��tIO�OL`�3��,3�!�>X �P�v��> ��r�@'l}!�+n�h��%Lz��Ձ3��y�!��-`{J��� C?N�\ݲ��7'�!�$*.�Xy��� �/��TS3��h�!�DQ�!��y�"�8�8I e׫e�!���.�E�ǟn�MrS�Zi�!򤔝=|1���+�IP�
]u�!�$@/̎�(m64�K�
7�!�pM���Q��X�T���7�!�DM�^�\=��䖃u偐�Ƥ0�!�Նin"i3��X��R��6�!�:�J��W��?}�}P�Y�:�!�D�%ei�|�1�	nϼ�rS�A2�!��<�4�٣�	LǌY�d �9!�!��7*��g��T��1��:?H!�$�X��
ƌƭ3������%+�!�$���t��u�Pjw�a!�D�=��q�'OC)m"�,�ƅ��^a!��΍�v�jpe!'`p!N�~B��w�h{wg�)#� ��S.^�дˁ���W7�3pH	������%\O�<Q���x�pm�ѣ̳-�R(���%�E�6]��=�f)�i"6�ɽ~���3Ee,5�@�9�oْєB�I#+P���/UYv�HTR�V����<]��ȳ��P����㤁;�6�S�\�b�hEeã/�¤;%#<FwxB�I8.P$�:�m�t�4G�l��Mҍ�
am�c�n�⠎M�IKK�08��r� �,]A�CNժFZL���s�@�ђ�9���;�KU�m*�͚�	ۗ	�z��G��s8T�ڢ�׼�p=!7,[��2t�d	��[Պp��x�'�2%�T%S�	�H�Q�q��!۴$R��HJO`���fU�DE����'�^d�ea[�+XB$U���-y�'�j\�*و��y�e��2���t�π ����!CN�������\�a"O1�S���BHp�0�%۱�}�!�E"�4'�p0ǉJ�]�')qO"tcs���r��X�-[4F�|J��'��-�ԅݙgl����k�/�$)�δ%JԱy���o9V�0�[�R�j���O=|l��W E�Y/���d�R1g�Q�����Ν?�P%�����.q�_<��AIR^�(1��`���+6"O�U���n����A!:V� ��O0u��aT8G�
�#���z�H�EKW�O��z��͗ l(�����2�@-��'f�0hQ�Թ2H� Ɇc�z�X4�g��V5L�)���Lx�����U��	��'�(h9R�B�"ItR�K6(�j
�j�������r��,qCW�o�\ ̐�0�f�+��"Q�t���I�%@�z⁚
�<}ReC6NC�OX�O(ɠ��ۗ`�6e�u�4x��≊<
]Pp��J�?_D���,�kw�a�	�'�`�c�H�!�la2���g.a�'ڌi�e�	��9�ta#%0�H��8ʧ��xdO�BRJ�0[���H9x�h�)B�z\v9���U%�������f"ը�i��
��U���\���~ܓ��<3ҀѼ�V�p��\������	�C+��;�h�U�d�B@����Ue��W�6�R�GF�l� u;�_�p=�TGν=��T�a�ֆ<���
h�'5d��qNG\Fjl�7���:,`��ش{�m6jJ����3��R�f��`��'I������.�0I��D�. T��'w u�Mh�Rtk�Z�d_�@P�t�O�|d f�̬�n 2�Ǆrd��j
�'�dŚ6�84�L1{B���$M���BF�)�p�A!�i��s��١P��'s�qO�б�R�<�D�)R��3/:����'=�ěDD�
P�h�JV�U����OQ�<�|���F�$�l`RU�ԝ����$MNE���� ��\���ܟ�Q�`���\�KH^	��5L�H��".}�8\�W�#�4�RqH��X��U)>D�8�uc�X�kb�Qh� pj��>D��F��d����#aP6'�H�;D����	��D�HQ\�ę���'2-!���@���@UHF)}m0��Tɘ�,!�$�Q��`�
�}�|��Rm !�$�:3�e�1}ǌ\�RC�;8!�$��<��U��>N��i�B5$!��&*r�J�!P�����q�
qf!��5�ݛ"NԌ��A��T+!�D�1b_���� ��l���mG!�D#k���s@��XW0���B
z�!�d�0Ν;e���:U�-CV.�+N�!򤄥r<d������>N�L�⭚%�!���8j"<�`k�7'S���fAu:!�DT&2�ڐ���Ǽ�e�&c �z�!��܌d��+�!_�[���s�B�}�!��/O�-XΌ�~P����<(!���$h�zte��d)�H��J&n!��Y<"
A�E+�+$��wꗍk!��M�gs��x�Y�kd�C��4�!���<\� �$�ڃN�d�S�
���!�$��F��0/[\�"����!�D�T�Ѳ��L��-�s��Y�!�]�)<��@d&�E�U
�n�T9!��&.�8$JP�[�v� �!a��_�!򴴭��_�2C���ZD];�'��鸕hϷ]��i^L��3
�'2(��W�.����gͻG=شQ�'�`��%6�2���͆�&�'�b��(Q+�R�6���dԕ�y-IbRj�ڑ/^%���μ�y�,^>_�<�b�p] Xh�+�y2J�3�KƱj��KbCC�&%����RTr���C�Ub��
x��	�ȓ ��Q�ӤIrT����1_�(��ȓ���ٵm��
!:� �#~�&<��t��舒,J�x���C�ܿQ�Dن�S�? �{u�۠���kA�LJ�sC"O@%#���%:p�9r�AހX��9��"O`xZç�=��*�*��@����"O�`�6�XM���p3���"O\�E �N���d"L-N8=:1"O�8��g�!�r��w��Jl̀a�"OZĺq��	Q7v�q&�N�iǼ���"O�8�uĊ$a��H�-T�/�|��"O� @R��$o���gÌ$f���( �UH�l	xX�h���S$S��ɧ�Ũ��՚��,D�\���!0����b*1>l�zF?D�����ljj��em]�,uHi�7�<D��Zqͩ0�Z+]3P�}���:D�s�łc�j��'<�褰Gk7D�\BFE�U! �S*D�k�<1+D�h�#*@-Dڼ% &GE<�r�)D�l�WN�(V>0b�GV�EP��Y �;D�x��-��|�蠊j������:D�(�F(�U��(1��+ *.]0*:D��y%FZ�|XQ#�Jc��c!�7D��(WMS� ���Q.
�-�����!7D�P�$GC�5j��
a5~�Bi!D�ha�7o89wa��vNNm3�:D��A%.��E>q�֡F�~\!b��8D��e�R#wl�C2LÈXi"�Q� 6D�tC �� I<1ڇa��0A�P�'�8D���rM=I����T��R�(6D�@�iҢ��eJ��3/���3D��#��՟Ql$�[��[�P��	?D�HBu%^�[}h=��9?ޥ��@<D�����J<# ���o��후 ;D��C��+^m��C
,yx1`�O6D��hW	U �P���{DC2�'D��vA�>� 8t�����!��#D��Z�ꎱ���f�8������4D��x�;2��-&��O�B��vL3D�z��=e&�ΐ=1��=�g�1D�x[�M� 4X�HM�y�تGK/D��ť�$����KЗ$6�4C4�-D�ȈEbXO�nx�rb�70�P}p��+D�\�B�4=t�ڄD�!/�QaL,D�83�[� M��c�,)���o$D���(� '戹4��%b��e�?D��R�@�A7�E;�Q-؀���"D����C�ZT���h�;g|�D�v�>D�̺��@�u;�Α:.��c�=D�$	�o��O��9{E��5�l�)(D�0���!(��r���7h�MpR�!D�0�M�2PY"m�*Z5M閍�b,D��葤�� �TaB� +���ړ�(D��3�Lۗ�"��P|xuB�g'D����N´s����N�S9�I�B$D��CO�3j�Ba����,H��rE!D�D�Q"�w�>a1��u���t�>D�Z�E/T�8u��(�$t.$IZuo:D�vj���)p��W6^��;��#D��B%.��T-.�Y���L\�$ņ!D��0mԕKn���e��(ĺ����?D�PR�!զ�=c��0
��*B�=D����h�pAA�+��.�t�d�7D��µ-��1���0�[7�l:6�3D��a�N��V�1z��G:f�,QAb5D�ܙ$ٶ_�}���F5@����3�2D��C�:�"��)�f��n/D�� �8 �Ik�*Qs!�#ZB؉e"Ox�Be>;gFu����*=4�D"O0HѲ�L�5�A�wd��5T� �U"O�p�iQb�~<���lG�qx�"O4 0#y[��R�;Ѧ��"Or�c'���q5~ͨ&$��m�t��"O�=��$E)a	�k�#�  ���0�"OJ��c�
K���B�;lv�8#"Op$�	��pF8�p�X[�Y��"O`�z�ט3��ٓB���8�r"Ol�q� �����˄C���&�#C"O(�6�-���BM�Dx��"O�A�ҙA�p�S&�J�2���"Ox=��ڰ$x���-��!�"O�Y�LC-Lw��A�Ss�"O�\ ��2Lu�0�-�	 �"O2,�#�):}�x��m��X8��"O�(@EY����f�?�99�"O�\�E�G/	L�#�Y�t 
� #"O����D�x�б���O�9c"O��Wo�)%��*�� �5��"O��tE�����*aiX�k�4p�"O�]��H�T)@����Y�"O�� ��X0��`�%G��T����T"O>3�,��a\���ve�W�`H�"O|9*�kԓn{���3E	*wB"���"OZ�81J�o���!e��R3L�ʐ"O��Ռ�hPũ���2�2�Iw"O�pC ��w;^�Ԍ��\���*"Ox�1�jS.�x�_�k�����"O�@�K@$^�2iI��H�T+؁�"OxT��D�JB��ƍ٤D#|D�"O����"}) �!w�@�b�,��"O�+�nL�d�h�8J�I��-�b"O�q:��ϒ9����&U�	��-�6"O��0��9����fF�Q�P���"O��``�n�B�	p�8�Y�"O�y��hFF湣��ڰ�n�c�"Oh�HIPT��e)Zq�~�!"O�}���6��H����C�"O���� tZ�0a��ͬv��""O^�3q��	����ϲm��A#"Ov���B����iQ�V�[n�=�"Onx��߳i�t�̅F]<	�f"Of���d��� H#DǇ7�*�5"OBm�W�K���M�t�Z=_�d�0"O�q3�/@A�<��`c���,�y�h�d@��V���bC@����	�yR�ͩ~��1�!US�C��>�y�k��L^L1���C|�t��A(�yb푙/{d���mǄl��pщ֨�y©&gb��X%K�T
�*@�^+�yU�K�buX�	�*N<B��ҡI�y"�L9xx�IQ���A^n�h�lF	�yRض&������3@K�L�3�S-�yBϒ��h� ��2������y2D�)�T�u�.B�F01Ħ��y2N�7�,�`#�##Sz���f���yb@_�&�s�ι �i�i<�y�	�[ATY��[�eb��:$����yR�
DL,��S
�;^�ԁ)a^9�y�C��J���qsز�|�TÐ2�yBT It8����X�(�J����y�V��T����� x�,(��!ڪ�y
� �j�e�OD�K���/��$��"O܍c��g��u�T�Y�Q��̘�"O䐠��"�ca)2����3"O�5:%�]�.�	����B��{T"O��Ys!� Z2��3/��4�,)�"O�����)-�q�.F I�v�Z�"O`u���¯h�<\�n� o�d�0"O�;�@=Aۢn��U\y7"O��h�eҠ��Ңզf^>�A�"O�h(��j���0ߣR[V��"O���-̦�	���JL�̐�"O�4�0	j�  a����D6�T"O,p����:}J\!�mM(NS�]0�"O�� ",�
5�`��]�i[� T"O`�5&�Y`�`0�0
!~� C"OT��PaF19�鋀 T�>�1��"O��C� U��4�0fS�K�Ț�"O&D)$n]�VR$<pe�HeE8Ȁ�"OҤa&��!���ʷ�4'^�i "O�(�̆��d���74Eb�Ӳ"O܍���N/(��@��l��n.�4�'"O6d��Ř�{F��E��DØISb"O�\#�0p��c�����p"Oj�)e'�p�j���q���F"O��+�A�?2	0L�v?D�di�1"O(���P�qy��8��I�|�,�#�"O� c�kB�#�����̮eB�6"OF@9L�5��Q(�$M^�M"O�p���<E��ڰፃ[[��AD"O.Hʣ��8RY�왆!OJU��x�"OP��a�RB=(� Р��� 4��"O��-��Q�d!"�ҤE*���"Oh}���*H.��'��!e�hy�"OY��"^�Zԩ��S�	nq�"OfE���
b���D�=
�HAp"O~Q@Wa� Q4@��
{�'"O�1#��Jx���&L��	��- "O�����7ي�y"���$��"OxѠG��L�����0�i�"O֘��70f�QfI͞|�x���"O��v �/k8e���#+�di�"OL��`�ӌ�ș�j�0���� "O8�KUk�+RL.v�z���"O�ᚲ�4"������s�n%�"O�L�D��A�1x2LE���b�"OҤ��g4T��T��C\h���"O��봮c
����[�SKn(�"O�1�S��%$i脩�� EEꌛ�"O>$���*8���M6l-�q+�"O(�3a%K�U��Q����4z�"O%�#l�
b"jm�e��.L�"OpH��*%�����7���y"Û���� V�L�3N �
����y�N��A�x�����$YU��z�m��yR��0M�*�N��F���F�L��y�R ����H)7�Y�O��y"���1�Z�㪛/*�vHՏ�y�ѻ�J�)�
Y3��y�@?Z�Л�Oޏo3f�S����y���'��3�揽�n �S$���y2F^�i�J���6��0���l�<9"�wH���e��H'��Kk�<1�8��}�rS��x� e�d�<Ѣ&C8g#����dT�`%�x�Q&DF�<� ��"jV�Ww*�Juşj�pԚ�"O�H1�l�
2��9��,�"(��"O�9���Q�~ ���	]Tȝ�"OB��'C3��ra�{�A�6"O$��g'Z>w2�ʸp,=��"O���r�ӢY�@ pS/�h�x1@4"O�4�FƢ�4t:q�W<�(xs"O8=����
�ջ3�I� �&h�"Oaہ�2�.��J��U���!g"O��cd�bl�);W`��7�4�"O�*L�yN��.5Gx�L;a"O�B"(ْ9���8<��;"O�$��.U
A�0�x��J#>�*�"OrTsb �  �   h   Ĵ���	��ZHJf)G�5u��(3��H��R�
O�ظ2a$?�K&��;۴%`�F#�M6&�ׂ�g�`y�C�%&B6m�禡b�4n������'����<��@b�\�ٞ��0�J�E�O�du�O���:��B�m��+@ �D���6��g!gy��H�]���݃����n#>�*����D�k0v���X��䘩 gE�Z,0����I<��ܟL;�! %�Db��sF�R*�ʓ+]�_��
p�VV3�u���m~2d#`�s����g�S���'�rq"�(:P`�dFB;#�HL�O�Q"v���(O2�YH>��%�?�6!�խ%s�d������<�'�,� �z"<1 `56|`xH��UU%����%GR�����3uh�I!�V���c�'5��=�Ci@�J��'��ADx��Bܓ�������L1���3#�Fyp�l�-������	4qH�� �/I* [�3�݈Er�xEC/�I#6���i4��P��Y�KN���^��$�Տ�<��<uX�pb�I��H��"�LN����l�vd��3�IV����69F1�0)��xll �C���'�l�Dx�`Rr�	� ��E��I9L-�8�-û	Z@��0���Z�x�^�Ԛ�N��Bep�x"M�0-&l*���O�(1t�G�<�-
6��oZV��Y?Y��, ��,Pn��U%`p�M�1.љ*�P0/O��ە I�K�'{4Ћv�ɾ��8Q��H�L��2f$a���6#����f��bɦq$��Sӌ��bԔc�ăca;���i�J߃)�D�ݯ9�v��;�fy  @�?���Y��O���d�� ��6.�t�Ջ+0 �0P�Bi4��ē��mM�T�O�|z��lz=�W�'�r�'�R�'�P�2u ie]P�ka�B�Y&�'<B�'�N��!_���	�E������
��&��'B�Y���R�5��q��� �'�'��/V��Mk�'�-�,Np�xgI��sl���ѮN�uўD��>L[�T���:f���"[-��듶y��1	,���H��v	�v��I�E�JqKr}�� �O>���O��$�O�˓�?y*���]Od�5P��1/6���?q�&�dQ��9�޴m ��	|ӌ�D���Y�޴,!�VO}ӆ���3h�ܻi:2���Q6!�:)ov�=���0r���D�z�� �W)V�wܒ �Wa/F�lAgHU0u�ҀnZ �M�i$��՟�i��ۄm̔TR��!���� ^9/�d�3׼i��]+d�9t� �g S�sn�E��ؽ@�Zc�!`�<en�!�M�w C,����HT8'�p���@jAr`	o,8��\9��6�a��l���mrT���S�d,yp�H81
�( ؍�C�S�GvF}`7%إ#���"��286:5qܴ{���hӬE9�nK�!�<p�;D��I�E�(M�T���bU, ) Љ��
�܌n��u�Tl��n>:���i!*�	Q4`	��^�� ڀ�	�1N�ёJ�.y�e�����'���'��=قuӶ�d�OXyR�"��?+��"֊Ɔ|�h�@���O����9D�p�$�O��S[�f>�aa�P����`��]�4�����E{�=O�h#ܴ.(���1�/��$���b�Y��F���6���@�axRc�
�?Q���DB=t>��r����0�� � ��'�b���Q��� �\#�<�	b���h�^���#�l�8r�� �+Գh5���q��O�D���&�'�y%F	������ ��V�Ԝ�y��2�d()�C���)��2�y� X�N��H���z����s� �y�A�LdFz�d@^ �s��y��=�j�@��7�����+
�y��(�q��*5)��+#�
�?yՀ�~���������(���J�f����$�(D��oئ18(�B��`%Y�D'D���f/i
�c`H֨b�0a� D�h��Խt��za��<q~��F$D���W*E���a5��MӚ��׌6D� �C	C��}�F��f�a�ɿ<q��g8�$g�������%%gI.9�H1D���$%��y*�H�e��3�*�X�C*D�D�RB�G�ݛÃ�0��� p	(D����G�0,���)A�d����%&D���D�6��w&�; �n�hϓھ�����V&3�4���d�!sYb�2%e� #ax����L�jM09�(���]��|f��|%�|�U!�"پd�����@YT-Ey�@	EQ�0F畺2�r��L#s+�cdlE>\��D�	���A����8g���Dy��H��?�d�i!l7��O�yRꌻ�
xH�Bэ4*�8ѫ�O����O|�d�ON��:c�PsP����>�*S��|Z�e�$1�O��	,8N��p��%'�L������d;�	¦z�(6��O��ݨ'|qa2aB�g4 7a-{B�I�k+�,�@[�.��]�'�Y#�B�I�Ul
	�g���ʐ	BD�V4�C�	/K%��ф�O�2(�2�;R��C䉶�]/�Jl�#�C�4���"O:̉#��k����.Ĵ8ՠe!��c�l��On�dͳ�th$��O���O����b�h%��K�9���l>U��a�FJ���""@ɦ���f�?_�zP�Oo��xsdΗ$�bU0u���)+ Ź��?v���sB�z���A$��+2�c>c�d��h��Ե7o��3n�܉ ��O�@�'�ʸ��bY����'��tg7o�nY�>}�x�@֯��"O: @Wf#'�~Y�bN��\���X�� �4���|�O��$\�E�!L�z��	��T�ht+2�I")�:�)��W����d�I�?���쟈�'�ҡ�aL7Y �`�G J0=����&��Ȣ�@?Ohp���kмZ����pc[H�I��[
Ɯ�N�����	�z!��q�����4�ME��L4��4L$ɔ��'oS8iB�yp0�'����~�'`�Pp��-�x�i�*x�
�'j�hV��.?�*�p�咹f��H�I>�u�i�BR�d�i�,��i�O���ANNjٜ�	��?!(���#G�O��DO�L�$�Ot�S�]��<��&1ePe� �Jҟ� ^�S��4�r�9 �"�����'p�u fm��/9P�醂;��_�4���P����Y��ӳ�0<��OD��H�If~�љhrl���@9�j8�����0>��M�U�X�`���@���p��a���a��`b`����19���	�JPN ��Ixy��/F?r�'��_>5�m������)�+>L>�r1��*m �dȟ8�	,?���s�Vk���L��
�ߟ4�'9���[�+��`G=}t:<Ir�=?Y2��M���I��ˢ	�Eb��
:��r���)�<����e�!ZdLûb'�"ѝ��[���O*��=�'�y��s��}Z��M�^Tb�P� �yb���<��8�$�Z<,�L<B�'�:��OiD�t��/WzH�!d�K��A���I6�V�'R�'n��grT��'[��'���^�|�BC��=1����_�1OTY�R�''"�#�J:|���i�%���f z�y�����0=q�����w�q7��i��[̓r3����T��Sɛ�Js�2��Pl�zsG$D����T��e{�I��+D�h�	��HO�I/��ZT�}�G��jc���"ڿ'S�A{` L  G<���O����O�y�;�?�����$IO�_�f��	�L��x�jF�f�hw�J-� -��L�� ��yRn��,��T�&�!z�s��M�~2�IÙ 
R�����0=��ጔ����Ej�Jd�կ��N>���ٟT%����۟�?1�a��8���I�l�;|N ���С�y���&R\�usU��VW$I���X��)����'A剴;�DI�O ���P�"D�Q�@�k혠�ʆS=��$�O"����Ov��`>U�"��t�\|%�� ƤULH
	9I�3jS�5�q�:O
�{!�D�H�r�O�uqۙV�DBC�ւ-���SB�'�̴���?���?WKɐG��T��^%�m �b����OZ㟢|���9+�i��H0{��M;�l�R���B�{�(�Xd�G�lC<(�g- JX���PyR#Ũ9��ꓵ?)/�@!3�
�O|�b�唘.�4qKW�ߐQ�r�"�n�O��Dѣ@��d�7[�g#U���'����8E���h�C�
վ}�a�_8S��I,!IN���&��I�5s4.]B�O� )� �BQ��Kg���
g�[~ŏ��?!��?9������ׅA�]��E`�T��\��&�|��'�azr]A�f�
P]�R�f�Z��V9��O�\Dz�ك	�hq���Ly8�2gA
�F%beɘvJ�O�剟\
�`�r�އy���۲��"H#D�@�P�
Ax(xq��K)��9p�+D� A7���!_j�j��M����-D�ē�
Du����V$`E�A�B*D�X��*[�O��Paψ�m=�*��#D��nT�o�fT��,�a��1˓�<a��M8�*��!Gb���ǒPh؁ f D�@7�[�L`p0aQJl��[E�=D�8#��O'U���p�\�8dTQ�4�1D�\I�MU�A{�Ԓ7�M6(��%yDf3D���%&還�ю�0
5+�#�O����O�5��Q�&�V��E�5ZgRA��"O�����*ID�Q#�	�\?�<�g"O���H�)i���7��r.�ЃF"O��ӣď�{�5m:���P"Oph�u,���8��Pc[�%��"O�	`!��@Y��3�a�)zr����I���~�r�D�b.^�c�ŋ
D<�y��k�<��	���{��y�!��f�<��ԌV�e�Rk�?x1Ne	 ,a�<ɀ�Ɩ)�aK�I�����p�f^b�<�Ǡ"l�`�ʠD�1Iq�L���H�<�4��;8�r٨�IQ�z� �c�KO��@x��(�S�O�d9���#��%��X��B"O�lk�J�CʒLb�oW<`���BT"O2ȣ�S�Ba��-8:T:d"O ,�!��}�����uS�"O�#�*lE�x��ڇ���!"O����ē	n��a$�J�<�2l��_�D*�i.�Oj�Ɂ��|��8q6"R2?vdJ "O� ��Y�.k~!9�̙wQ�
�"O�mr����3)TŨV@��#�"M�"O]���) Jh�H4/�}�<��"OH=�
[�dCRx��W�-p�s��'�f���'�>x��ۊN�F���N-��a	�'��9�E�b_^� �C݀Wݸ`��'C�E�ɌDv80��GU&@�L���'o��X�����$��nO�C��հ�'$��R)�Y�� ���(7�f�{�'�h�pd/��t����7�Ѹ(-�X3��$��e�Q?��E
+>���kn)<�rk��$D�|�dL�6����E�P�,8�`-D����˞%	B�3��O�3��0٠�6D�����cPDIqa��W���6D�<0�Dba֋I�7�x�����Ox�B�I�jS�8�l��L�N�j��ܕXg��d�?l6�"~��]�O^~9��1PNM0�	֞�yR��3p���Q�� �L:fA2� �y������)��VC)���'>�yRc_8|����*@��e�&���y�آYb��UL,!���2u�A�yҁ�C(���P�"��CWcŊ��$����|JC�B٪�hϦ��̂G��0��[�N2�
ݰZp�4�Z7G@��������MV�_^���2o��.8�݆ȓ$��1�֓;�t����/��m��.�`Q)c�ںfv������mvn�������ɻ���G�J�$��<Xv�VRB��9>�И���M�x�ִ� �
.]�C�	�ZM�4±IY;-7\I	����g>�C�	�>�č A�ŢW���"��,��C�ɦZq���D���{���`%�	�x C��!M�n��BkNt��])�%C:}��=����K�O�t
� f,hB�,q�����'���YR� )�<��a�n���'������	��@8q�T<^� �K�'^:�+�ʄ3�D�Q %�e�~��	�'��P�d��.S_V��J��T�~=��'��Q�G���i���GԂ=�>���Ex��iлI�� 7�9��E�R-�B�ɍ>�֜
G��y+H�JEA�SnJC䉱a�������.�7�L*iZC�Ie�`���ٚE/J�X4	 c{�B�ɇ��`�6�X7Iޭ�$J-I�B�I�P®��p��gqƵ!gH��k5<˓G`8��	�n��uⳎ�0���ӃB�Ob,C䉰-` %
D䐙h�4�Ѕ��*C�uP�p�4��%r�Z9"���w�B�	67�����j�l�*���T�LG�B�	.XfU#'C�5^ì�ʦᑤL ���N3��D��n��D�B�	p���	<o�!�d�2'��P��SBT �P#P� �!�Ѥpo��K��^�(���7�!򤒗�8�z��S+8��X����!�ή#�����@�9zz�4)1)�j�!�#e焸Ǭ�8i�h�3e$wў �4�&�'��S�ݳr��xy��k�����*��5���( ��M
4k��ɇ�Q�>���]|.�	ñ.�0U����(���`%���AAF�(A�ȓ'�:�"����s,6�X�}Js"O�$���16��X�lءs��}���'Tᘌ��ӻ
F 0 �Ö�J��R,�p��&���;�A�Gf,��
ԾV��X��S�? ƴ���?5��\���,��u�p"O$��W��Mh�JL��:�J<K�"O� �� ����P7k�,�h��"Oy#¢��g��ؓs�A�(Ղ�ےR��ɔ�1�OΤ�f��� ��Gʎ��"O���ՇʶC,p!�z̋T*O ӡ�U�	�P�G��VT(�	�'0�	s�`��5c�tIG��:��Y��'�<��!��/I
X�F`�!,tn]B�S�����a@�@�*�"a��1�V-��8۸$�B�\,�#)��"	�9�ȓ<|	s�c�4_����N���ȓT���C�� 9O0U�!I�)"��i�ȓ	�� $	�X���M�(����F����Û�Uܘ�6 ��؅G{�a�֨�������q�l�a(��&p�"Od�`��ro4� @�E�pm�ِ"Opa��9��%8B)?|UB�"O6�ӌ����ū�-�i7���#"O���g�I6BvD`L؞m}����"O�9�hfP!�vAGu�1�'p������#mOF�ȣ�I�J��(hR盜/h�����iV �:I{b�2;��B��;(���k�u��`[ 3
��B�I�9Cf\Z k�=s���e靰-fB�	��r�{��[PNȹ���I`VB��7nS务��'��8��n�'�Lʓ4`����# U��Ń�';	+Ԃ׎_�"B�	3&�`�3�߄m���j��(�@C�I�(;�;���.!Iƴ���ߏ9��C�I�Kj@��	B�[�^��n����C�
�r���O%l�y�#W�c1���Ĉ8����;M$���-,TĶ���ы�!� ��r|1�O^�kV2��v��Y�!���3^�v��ѥL*!�� c���!�DĈ"�<m�#�Ƶ8�$<z��Q�~T!�dZ���9��n�V�\,s"��qr!�
�� Ց�e����@�pK;E�ўP��:�C�V�����P(�en+�@C�	=1gH ���7k��ЪW#Hu�C�	�'�L1ॆ�_���Q$d�w��C�Ʌ1�����Ή@���rDI"R�C䉾qT��q0�@�vl�`[���3�HC�I��)1wIW�Q.��7��^��dD�h�"~�(N?KÒ`�rÐt
��R쓘�ynoԾ9�&�H�7<4 �Ż�y�e׿#"80��m�2���Ufф�y"D]O!,(���X8Nb���̐��yB�<9����I�f��d$R+�y�(ȮS�:)q�B�\�Jh;$����$�>o�|�!�NK���a�C���a��V��y�+Z� �i0iX�h�|��"!��y",�êUۂF�1d�r�9�y���d���0����a�)�(�y���Fk��a ��
��#CΣ��>1Ԭ\?��ȐV�$)��GI�X͜�I�J�<�6� �Đ���.&���JE�<	W �*vw���.�}�\d��eH�<��I�q�v�FJF�$�V��e�C�<Y1���j�5��O�V^¥��|�<	5d�f,\ #�\��x�!g\B�'����iCJ
���a��&\��I+A.2�!�dA�BT�����2xp=�����!�dD-J1�q�ͻsl*Z��=�!�� �Tk���'%%e ��y뤝�"O^4�V-�$�pQH�$�N͘4XT"O�LX�!���=��@Y/b^���'�|�����yR5����8�E��N+ I��X2&�C���}F�R�}d>`�ȓ��=A���B��� ��S!h��ȓ8Ѡ�:�[4w $��ߨ#�Ԩ�'-�qG,=:9d� ��E!"6�uS�'�~���l'?�v�Ka䅼b��+OA ��'�ʕ��$� ��q�3=��1�'9�A�#	�Ve�%��\�m�%��'��<A%ܠb����c�q`���'����I���Ɯ�D�@;z�'RT��cI�<��u!�I��p"> ������j��7"@=��)���/�̅ȓ8z�[�C^�s2ڽy��6Z`���p�g��TN�A+�d_.��g��'%�>�Rŉk�hM��
�^�H�!�7k'F�j�BG�$()��o������!�dR������E{2��˨� ��)�!��@y���;��"O�S�)>������ST��Y�"O�]�'�՚hl$U!G���,���A"O�L���i�tȂ��\�_ò�*"O, Jŧ�O�`,���Q�TLJQh�"O�h��	2H�D�8JL�H4r3�'�b�x���S�!��щ�e�5 B2��G�����>�rW�;Z{� ��2�v0��.���&��%b�v&݇E�.E�ȓ,��HqF�B�P����]JN�E�ȓD��1���HȖ}�Gڻkj���Ɠ1P�[��8����(Q1 �@hȋ{��ؐ��$F<vy��'�ҙO9�TB�#� vfbm{�M�
$.�8��^&\����?A��"i0����I "Y�2k�>ͧY��T �HȅU�y������D|2N]>Oĉ��X�>���t����T��š�C� [\Q�2��/R����Ob>�� $�p֎���.��gD�<	���=)Ć@l����.��5�����I��)Ĳx����{�����R��9��Iޟh��O��R%e�
	簥b��Ф2GDy�3O61���16���Ba��o}��I�#�.�۳�]�J��C�L��"<������.M�2�,է��Nu%��<	f�P�gʁ(���0�;O ����'Or����f�~�	X�j�xe��Y!��$T�ȓ���Pc�nݪ��鉴!��eF{b�9�'u�"l�����N�j�'�]��Բ���?a��E�^J"O�-�?����?������)48{PO��c�|swL@�������Ω0�TՉ���V&.����̟f��>IAr���҈D�#&��d��'�ٗD�(�6`�$õ+O�8`�?ѱ�4�M�R�������L�:�)Sc1)���K��*?ic��֟���Y�'d�½h���s�T�qF2��¢��mD!���!X���פX0Ѻ�ȑa�=�"��|b����D���r	�@��&%�#H�"6��y� �OC(�	ҟP�	؟���Ɵ`�	�|��W�v�RԙvmQ��Q�Ūs޺	��Z�&V܇f���B�	s��h�4K� q&́z�)�n\Tr����D�fP�A���6ǅ>�Mش��O�H�'������3S����X�f�"��'�ў�F|r�J�}�t�$ ��v��k���y�΄�t�z��AoI"E>i�fD�'���¦-��pyb�5��'�?�O@`�X��8X�|�٤�ٔZ�:����ob�����?���t�D���0i�<���e��]��Ou�5�'�ٰ�fM�$ y��ȉ�Ą�?��g$Ф-��4�é�|�� ^MJiq[��:��I)w�h">�4�����	Q̧��y��Z*Bm����9����'z��'A��h��#X���z"�թHlJ���7��C����^ s�V��g�M*���q��YK��io��'���78J��	ퟠ
���=��9�q-H�)q�	�'�㟘CïԹ-�������gb�3�S���\#T�t��c��9:����F.��$�,6W���rfO ~ٴ �"0��W���F�����Ǒ��� ͓]�`������'��� ��P���-��d� ��pW����"O� 8�%�9���"��Z(@3Q�"�ȟ�(���#@v��#M���vQK��O���O��A&�I�=����Oj�$�OrU���?���6v�	�"�W?d&v��aN]�D�d�'Q�=:��J�*��� ˟�h���4�8Z�柸9����>h`��I7t 9��\9�@�g�'�h��C��[Br��`��u=B��O��*��'�b�'��O&�S �u���L/ (ЛU�t�,B�Xdh��aŵTfNqc� A� �2�d	S�����'��	�2$���AcH �ࠌ>3C��F�
_4��I�����x�SٟD�I�|B���-f�P-x�B��%p��'Je��(�'	�t���ՙxڷ�I�=*)�	ȯ	�$L�YE��Ǭ�0sִ��<I2F�P䉞3�M;ݴ��O@�kp�'E�IH"�_�V�����m*`½�G�'ў@D|R ��X8� �&`s�됡���yB�`�Q/b&�"���S��'2\7m�O ʓy~��ܘOI� dK�p�,�a��}����DC8*sh�QV�Ԛ6���S�K�!X��0�(����En���F�p�o�BG>9S�򄙩�r"I�+��q�k�{ ��R�KZ*+�J\�C.N�l���,�AGz���1��'���'D�鏻i�8;Ug�2���Bbi�l=��'A��'��R>�ExR)�af��q& .��S��+��>Y�]�x��k�GwnD���2-7�K�
�<���ߛ6�'�1��X�`��hQ ݹ�dT�ɾ�	T��~�	T�'��,p�	̵3/2Mz0L�5nr����iU�'�&5�|��	��j�������<Zv ��CHG~b����7}*��$C�N�T쫃�F�9i(�9c��;EL�q�!?�s�>!���Y�$�x�Ӵ&���"!�(פu0��
2|�]cR�>�p�O�}�4�B�2 �/1��<Zf���i?�ʕ	Do�dTq��K� A�t�S�e�@����7Sș�a��'�������wCEE�"Y��Vi��y��-`��1$e�oԆ��I9��I)V9�'�z7풳�~	�悗P�d����X�I�_��'�,#��hG���qb�Ù;�&1��ϑ;b�dM��S��'d����O �R'E�g7��ZA�=���;�c��uR`� �@��'�j���'C1��i���!�r��$�F�|����q�'����8����9O�y���O q@1�P�W
��3&AϠx�(�*��'Vi���/z�Ny �G�i=6XwCH^��C�ɝ��=
%�ްOt,h��j��&��7��O2�O�1�����|n�Q�leY6�5,�x�g�JT:��䓺hO��r��r�)��=q�턅t�.C䉀��h	Q��<v��i;0oğpC�	-uɘk3(�)+9���u!AK��B�ɿp�*E��-,_dȋcg���B�/G2F!A������@O�d�&B�	-l�,#��ޱH��i���ʬK,C���)��%�Ir��D�ȯXK C�I�=���«ٮB3|U����=�:C�	:�$�����U�X)Q��<�HC�Bxe�$t������ؒ�2C�	�_l�I�g��-�p��\>�C�I��S��ۿ�c�-�_�C��=`ޮ�+Q��z�6�)6������2��аxǬy��" k�:)c�()�4}k�M�2f�)���n�`�)*X(|)�Ý8x��ƈĘ(�Z5���?JE�,h@��Z��<�-W6@ȉC���Ik�a�!�Of� �h�&]jT�u��+z�0�	��u!�)f4R����7(�lQJ>���$i2���B��bO�R�FC��>��p�BoD�(�B�;&��?~ C�	3ˆ�@�yj"5��"�\C�B�I�?wش�+˯i�	��G��$��B�I1e�,Yp��R�4��C��,2ZB��6^�
x+a Y8@�`'��<�,B�	*.��x��鎑PH.��g�B�
XC�I�!ZJ�hsIA�&��KxC�	�B�ڠ��<��e8kH��jC�v��9sҍN̊u�s��	j\~C�ɦMC����+�8��E�[�HC䉿e�4��q$B/4zIt�D�@C䉻JD�+�*ϪQc�xt�ߎl?0C�)� |�j7�\.�qU#�'� %� "OB� AB9�y����jM��"OpAe�/	�y(ACN*N=��R"O\��w��]NЉGA�Y P�z�"O�D�4%O�A�ZP���N	<�PW"O�iJ�G@�FnT԰���3V<�P"O�,�b��h�T=���?"�����"O��b��8�.�bc߳8W`�g"O��ǭ(ղe0��ۈ ����6"OLA�7d�&m~�QBM�V�R=G"O&8��,R���I.
�5��"O����L�%�|x�6'��f��<�5"O�T��ހ|�����Ky�ĉ�"Ol���ȓY�L����S�.�4�"OvA�T�g�PcIݸa� B�"O~�I� �0Lz�ȵ╭KЌDu"O�hwe�b���2�x��f"OR�&Ѩ-2V� �ȥ1�ti�a"OT��V�06���!��.L���"O��{��ѠDri``��:�d\	�"OB���%:$�\y`֏��f����"O�l��M§�B@�T ��#��L'"OT���5%V�rPn��Y}6�X�"O��bzI*��(u����e"O
mArF�+<��Bb�#oh��"O>�q��Xy�����I	uh(r"O��@�����JH�^x�!u"O� s��5"���C,P)��#�"Oֹr�ʗ�Q����� �B�&<+"O4�1��sL�31` �Z:v1�r"O00;5(ޕ���@�/;4�0�0"O�|!�又}�<`��$��.�t���"O��p'յQtɠv�GK��li�"O��el��m��MЃ��+�|��3"O2���A�|v&X�B��My�iW"O��a��=�Z������<вp"On���@1����ք�V���"Ov�;�˕2ςM�1��`�(�A�"O´qB$)%��A���Y�	 �`@D"O�9)u�_������@8ؔ��"Ov��"K	�8q�U��u/��C�"O�ш�,��E��Al�v�$�"O(����A�_}L��k1�4��"Oũt� !ɪ���_%���8�"OD0��5A�P�㊏<}���"O��2��$�6�H� vF ��"O@��T���趭�5t,�i$"O���e��UK�Z�iW�u��"O�8sL�	:1��?>,u�"O��Pt��-X<UR񲢺���@�L�<1R��jH���P��,�j$��&�s�<���QIr�HO�@Ǟh�Q�Z�<q%!�8F@\����nnRd�GL^o�<� HC����D$ϻ�"��B�<�QB�V1�lӒj�1C���:��S�<�E��]ꐜ2t�G�s2�P�<�2��m��e��@�5y��r�DE�<�oD�# �}�R� ({ ����<�E�V���	'�\#�Lw�<	�)Ε]�8�@�C��L_�#��t�<١��f���"!�!u�U��X�<��ʑ��u���s�z�TM�<�E <�L���̏R����I�<1��[8�B�2�/R�PI H^�<� �a�G_�hB�E�5�X�sT�|Y�"O��C�jL�G����&-G4Z�"O|�p�O\��,���>/T��"ON4��J�>j��HC$�)`�!�"O�a)AG>D�zw�L�u�"I�"O\y����E�2i�i�0�=�"O\�9�P<��v�L�=�@�"Oֵ�e��1	I|��B`��C�m �"O�hJe��*�!��͋�e%�B�"O��C�*B�[��1��~��:`"O��B�6��Ċc�ܰ\�,� "O��K]x9�J$�$|�4�"T"O���$�6�|pH��+����6"O�I���'��)�b���up,��"O�葶
��i�Z� �̞�6c��"O��HǍGC�b�У(��Je"O�ts3$�G��rʒy���"O�0�#��(nԩT�1'��(S$"O�9�:sQ� '��$ ,m�"O�ỷ��h8ii���Yڣ"O`�D��$c�(];��KB��"O|��@�d�֩[������u"OD�ذ��j��k-v舰X2"O,�곫A��M�P ˊԘ%	�"O\�jC��_:��s��Ǧ�r|�`"OD���-�E���.�_�5Y"O�M�T����,9��@�b�5�P"O��H��!,6��Cl��c�� �"O���"'�9k*�X���ؐ��EQ"O���HM��0����Y���P�"O���b�����7@��y�C"O�4��l��8P1/�'ⅉ�"OB��TDۊF�8��`����H�"O��s��ja�Q
Y �>H�!"O�����zמeI�nZ�?���SV"O�\����!HX�pCm�F���"O�).Ӟy4�k�.Rؑ�"OJ1�aZ�nx��쁮,��(;�"O�r6�� gJp�;�LB�r�sC"O>����ڰ=�2i@"���~�S"O6$����2���`��C�9��h��"O��C�
L:a�&�R�Eڕ`�����"O�X��F�)IMN0Z4F��"��D� "O	BoR�cA<�E�V{��q"O��A��Vs���ذfD4���"O`�	�??����"C�*h�!"O&�1�<m�<���BA�t�:�pU"O�J^-@��v^-G攀т"Oa�d�D�
��$'� x��"O8�A�lUf�h9d 8xЌ��"O�Q��O�C��P�sݤpQ�"OR�H���h$�5��cڙG�}��"O�+�녤c�n�pç�+z�*qaT"Op�A�CѺQ�"aK���F�j�3"O����$t�^�0�e�,u��=*�"OFL�F��3cs�!�g/��8h~�H�"O����%̮L !qN tp��E"O�S����@���`�\�S��ī"O���ú�a�qnO��=��"O,X��1Z����&�sܬӆ"O9 0JP:$�Ԩ����$gR���"O<A�q�Pv$ �U�F��[#"O��)1ϗ�4���(DA�B�Q`"Ot�(���z�e��ز^(��"O� ��`�q�<�s�R1%�2X9�"Oii��4=rE�0M� 9jN	��"O�ز"D��e��hu�Hqc���"O�<ȁ�T�]��FkW�\EJY#�"O�A �B�'�D��S>-1�H�'"O�Y�C�x������*�;�"O�遊��8YX�`�F�n
QBF"Oܘ�5��F�
a��$�FYpt�e"O�=��㊸+���3��{O!c"Or(AL	�A+D k��R�2��8�"O�I� 	Nt�h�š�b4(�"O�,��dΆG_�EZ#-��P���Z�"O$\�$(ۨph����"�!(��c�"O�4���J��Q����a�~Q��"O�1�(�!S��B�o��xl��ʂ"O�z��Ԅ��G��-&���"O�,��#u�Z C��';�q�S"OB���!�ՙӄL�6!^��"O���vmI�3�	�uJ�be"O�C�$���l��G��3�\�Y�"O�t�%/��r�@S�d�>z�D��"O:�#@�Ѝ�&���2e^�"O2�`F@�+\xe�&�ԕ%D��"O
|�`�a(�]��Ę7Y���"OZ0a� �;jX�\J���](@���"O��sr� *�I�$萗\#|i�"O���Kʹ%J���ˤHj|�@p"O�iٶ��|J �����N�̊�"O�=��6_�@�*���U���h"OҘ���H�Ig�(�!�*n��8 "Ot�HT,��G�R�`�T���36"OHE
CkB��HB��*"��"OLQCʃ$6팀�"�L�!�aK3"O Ց�N�E5Ԣ&L̂*�F�@�"O�çI�jI��1�TV���(s"O�4�%���g0����
/�>��"O�%Ǒ���|��N%��� �"O�XP%BI�b�^)��ŀ�i�,��r"O�ĸ�-��E�"��vjگ%6��"OH���ͯ�: 
�� ɜ0�H5D�tp��Ud�x'�]�zJ`H�4D����!:�R]9� m0�`�?D���/�Q�����ߌ�X�d�)D��*1�ݣN�D0rG�!M<Y�G)D�@h�)��C=L�z��;eh����(D�h�d�1h�]�0MX2"���A2D�l`��
5l>,B0�H����p 0D� �u
�d�RC�gF�z�����-D�,K�I�&��8�3�
I�`��*D�`�	��<���6���~&��A�;D��
¤�66�P������腐0�>D���"K��5'�E�A˝_�!��>D�4�$�ψf�DC���v��QRV�9D��#%��5���� �>e��P��:D�<X��\g��8[��B(��""=D�H{��K���b�_�K,�4y��9D�p�%GŕPp�hФ��2��H�@�:�I�^�T!V��>j.��QB�6%ր�O�͹�$U�3���T.=~���"O�d+�A�}�0$�D�#Ef4!�"O|Q{qm	7F�Ĩ�S�ʪ
E ]��"O�E��9���H���"O(1�2ˇl���r㓹va�� "O�}��"�s�����_3�Ѐw"O����� vS�m�p�H�@(3�"O� �D���C�6���A�6�-��"O>��2�F�#�[Saj�9J �X1""O<ځ
P����؁�³<߼U��"O��#׎�&Pg ��Ҁ���@"O����صRZ�a�T�L&vܠ�� "OFu�ҎÚ{#:%���Qlڄ��"O*��2c�)\�p+F�	�2t���"O0j5�':�؄Dh�e�V8�y",ٞWVrX��%A�H�๴n���y�Ș�aF3AO�y �4 ��J!�yR�C�T[@ej�.�oz�:��E��yr�W�U.(�� �;j9�pq���y�$�9A6&���C�T;������y��9��XK6g�/F�f�v�;�yd��\&U�O�4��i�o
�yR�K7],�ЁE�A�ym4�s#i���yr䚟&L25Xp��5uF�� �¬�y"�V��^�r�GDE�����&���y�O9�$m9楁=vO�A�D%֢�ybK��Qz%�V�v��1��I��y��φ+B�m�'��m�v�2����yB���_�f=�AjQ�h����nɧ�y�$� vP��1.ń8t�l2 ����y�`���ZhԀQ���aڀ���y"I�)j\b����a0W��`�C��"n,�A
gH*P�j8 1Ι�0�B�	:9( � �^77:@�r�.�B�IN�1Ѷ�.t%,��5S�d�B�	!H�� :���;T�X=�%��57��B�	QV(|�B�
nKrܑ0�[�<�B�I�:VV�� Ub���';8���m�j���`�.^�3`�`	�'����`F�a���c�_��d��'�,Ȱ��~"��׏�=�M1�'^8u{5m�#�9����L�l5q�'Vd�QłD�0��5DE*7(��
�'aTM��!A^~R�U�9�*��'���kq�N)�F�z���&%��"O�d�Cm��mV�����
c&f$HV"O����!}~0�çGK�c|0Hq"O$�e��2���9����N��Z�"O�y�W�A�����
�!�~��c"O4q��Lqo��#�i�jg�}��"O~�ط��;����T���S�ΜJ�"O>H�e��',I����V����"O͉���gh܅���$�gf8B�I�'sL0�!*�tQ���U��PC�IA���  ��J����O���B��.vu� h1U� ��.N�=�C䉹/��� ӯ_,4��%)!���C�#,��(�.��1Ȥh4�L3�C�	6;��I� ͯR����Q��.wjC��){��@��9-b)3̐7!*C��

E�X��b�5�����o݁uԴC�I�Pub�.HwM|�����C�I�
�\��� �x[<@h4�ҿE0�C��&w&|�Ă�4;4�"�(�RC䉉L	FH���U����R�^��C�I�%�v@s�	U�=Μ���:l�dB�I4��)b`���N����ɪ`��C�I�PB�A�kH��:A�A㖯P=FB�-#@�
u�IM$����;p<B�	�VNdP�t�	$t�.]* n�=B��|���h��P�TPJ��	�� B�)� ��9r�64ȸa{f��%Hċ�"O�M��-Ԋ:��lyp!ۺU�b�K "O�b�E�m��9���2ϖ���"O���ȺsZt���ͽ,de��"O>��AIM%��#SN�y��x�D"O�`�u�U¤�2�BB/wN����"O$�b@�<%'`5�w˿%����"OЌ�N�4 �.�R�M�/?,���"Ol &�L�Cz�jvm�Dc���"OJ�+���z�f ��4P�1��"O���P�s����3b�2��с"O$
�a��P���@���P��q"O(T�E���)�� �*U��Q�"O�9i�<��(����!�beB�"O�	6�/xm�c��+:��8"O����Q�nn��0%I>�JAps"O�lڣIׇFI�e8@�Z.��u��"O��سŔL�X��PlI:f90�"O��2�׊
>0��',F�H*I��"O�օG-����� Ė3�:�Z""O���*ɧ9Kڐb3Ac2��"�"O>kVfT�_謄�"��Q$��{�"O*� %N�D�p��zx`�"O��0��.!M�%��=)�R;�"O�����ҀK�L))�"ќqa"O�8��hɅN�|p(q L�H�AP"O(r!�Z=Q˜dxէ�=^�Y��"O����	���5`]�6��g"Op��ʢ.��hA����
y�Q�"O
Ik`ϥ\K���V�wR��"O����S11�D  ɍ�4z�Q�2"O~����d�V�Q�����j"OҤ��L �h�ɣ�ꑸ4�FMh�'~Yq7�6������WZ��Y�'O84� ��$$z��[�_<T���2
�'!^�j2�����аu�҉��'�RQ@T-ܣ�W=oF�`�'U�(uc@�za��DȚk�r�H�'N�;cKiNfa����e;p��'��尐AAj$����H��c�'����Âܑ]�T0��U/^��A�'�h�M�,~���X��73��X
�'cι�ZhĢ�J+y�h�ȳ���yB
m����&��m�S���y�N;4��Z�h(&��(3��.�y����H���!�&]��g���y��P8��e�G��Jt΋;)�,C�ɺpk�p�A�!#�`���-�:GBC剳=�\s2�ȨI����+|�!�䝜ph�#��àX�P� �j�@�!��B����46�=*��Nx�!򄂦S/�����<!:5qC�z�+�'Pcw
��R�6�Sb�8L4���
�'�Zͳ�C�s��r��&`��	�'q~�	��^2g2�Y�+:�Ќ!
�'�x 7ުz�<��0 E�<�@�K�'�``i��[�#CMB�CĐ53�%��'�����KL{ �{T�V�4�"!��'Q���*	�]���*��2
�'4�icsFC0z�>%���84� ���'�T(`��<*$���A2V����	�'Ϫ��ā\+y�Fh�`��Thت�'�PZ��D;T�A� m����
�'��0s�˓�2�a�'I�![?>��
��� ���Av0���j�%�"OB貤��XߠQ�a�ށ�r-�""O.8��"NA�y(��w�tJ"O��! O>��u"V�DU�5P�"O��Y�8� ���p���"O�a3脬�0��7M�"D
�"Ov5��W�j�lQ�rA�^��q��"O�\9�i�8j@�:ǭ�Q�0��u"O�IH��53��0⣂���d�w"O졲�IǓ��s"L�9�hh�"OR5��Ě%hʄ��A!`��|*%"OZHL��l�r�����"OeU ��.@Lx;S�ג5>����"O�����u"����N����;�"O�IKS���i���j�
��u"O�,����r���1�d�455z�3"O��sB���X��8��E�s>�b�"O�UӒi��nE��"!`�>
��{�"O�0 ��*	[��s�'�4��!w"O搑�hD�{�z��Qmضz����"O,<�F��714��ЬP���H�"O�ٰϔ�\`䝳�c
�O�^iK"O�×��,mh⍳��Z>���A"O�c �L&}�Tc�Ŗ
�2D+"O�DKSC��T�`k!G�։��"O�	#/�:$z�̨��%be�i"'"O2@P�è<A���ui��"Od�lR�N<�ēF�ݎo@����"O�����H�������@"O�=���ר_3�
��
{�����"Ob�j��

N@䩐=a!�{	�'�#ʙ=iK�IS��ĥP��
�'��횠�

Z�Ep0X�N~Ix�'��$Pf^'9(���| (���'��Ô�"xtl�'W-m�Z}�	�'��1�`��C���a�1]b�	�'L0�(���*�4g�;/йH�'O�����\)ab�F��v<��'��,��H&,I���L�5�L��'�� ����
������+���`	�'x�Y%%աJ�������{�f� �'�P�zjÈ)�i�Wo؄t���h�'��<�HM��r����f�B�k�'���	���8HDh(�p�A.`���	�'P��ĉG�"Nh������'Dn|y�)�:���VJ�{ �'o\(1����2��U@Ճdz�K�'=���@ ����������V���']JM��@�r��9�*�	9���
�'� ;��G3B깪0J՜y�D��'^z�������~AA�G 82`R�'���Q��-@���s���>+��(�'AD�5��b@��g*)t���B�'�E`�霼M�u�&I.�`A:�'��ds�k��i5����B���$tR
�'�TyР�D�j�ȧϚ�!LY�'r\��#��D����G�?�\1	�'p���V�J���@�2P��	�'�P���?|�>�� G1Ib5��'K�y����&hI� x��>.�0�'<VM��eF�fY��* G�^BŚ�{�����M�n�=sB5ʰ�_��a���z%�LENݨ1'��}b��ȓ��}�t�� ���Ŕt��p�ȓt�(1ا�ǖ1�� �.aL���S�? �@���+(�1��.eD�L�v"O��¥�n�Hm q-D�u+�X�"O��*ޓV�I���%_,��e"O,����*Irl)"c�I���b"O�}�siy.��GAy�\)�D"O�IJ�� o��Ɂ`���Y�\M��"O��#�ׄnX�#fG×�D��"O`i�fS#)��kƃIl�u"O �I��	�j�*��A�Iz���"O�;EI?R�U0�)�+�u��"OXD��Ivo���A)�y���U"OFQ���Th)"x-iz
��� Q��y��5.��Q�_�I:��c ��yR��6 �Z�R��I�n���S����yB�%�0���(�T��2E��y��a���@�&R	i���Y�yBDQ�q� �K��5Qcv ��y��ޤW*����i-W 9�c�8�y"�H��X�"&��LHDHZ2l���yI>\�d!囔U�P��.C��ybc֎��djg"�O�n���ԛ�y�ㇵV񎰃����Kj,e�vK�y�`A2Lw��YP���#�9s&��8�y�KK�EzZ������eb�8�y�͗��]8���	��'j̆�y"��y���a4�}>1H6# ��y�拞�حc�G�% S��;1�ۜ�y2d�:`%8���֊e��⟴�y �	�ejSB�E��{Q����y�������Wn����!1�i���y���E���7�X�j�Z��\��yrs>l�(Wg�--��ĵ�y�-���(�k�n׾����4�y��ȥb<�=���6aM�lh���yR ���b�14��Z�`�g+�B�,=�8��B�=�����,9\Z�C�	�l�]Zg���_l\�1��1W��C䉪K�&%Ô�:*���A�� b��B�	 p�t�cb=�*�����GؒB�
6���:�%��J�eK0F�PC��4GC�d E�-7�����[>C�I�!�
��H�*C��(��(HiC�ɛ( �Y!tK�~ъ���ӷC��B�I1 ����SN��B��S��0�C��1{�Ct�Q�?�2�0��9��C�ɽ�R��-@�KW$����>��C�f0��&O�3p9��Q�K��~C�2C���W�����FL��B䉖�u�V#�c+��5B�}��B�I2l$��2`��eמ1zЫĨJ�B�	9x�h	�lQ�sS�=��mD50"�B�0p�|����HO�y�uk�n��C䉢hb�+'$���ʉU�ϴ.TB�:����K�>��[e@�x�B�	<8(�����
�@ˈ��V$�J�C���&p���h6: �f,�6��C��1(���[ O*\L���lG$m�B�I�Mi1zu/Z�k��)��a��BC�<�2�j$�^�4�X5a�e��B�I�hX(���M)W��JGD�:�B�	�Y���C��2G��L�6(��V$�C�I�!~4�C7~�ð$7I��B�I%�]���K�-��4� �דY��B��n���$��R�6�I��ɜ��B�)� R� �M*%���"�gY	C3֬bf"O�t�����C�T�r&S�:,�YP�"OX- E��?v|���fοbN���"O
̸֭Ο��r�K��b�~�!�"O��cF�N
?��P��� �)s"OJ�p�k
J�ĺ�a }�4�B7"ON���i�6.��:j�'J{f�b"O���Ŕ�&�H�l��@��X6;D��� dƂ;��Ţ��6�%���7D���������a0�ΐMj�x��`3D��rł�r���͌E�P%+0D����+|E��A�B��al,D�hj� [�n�-ʆ��� �>U��5D��
�F�Bʜ�#�-6aA.D���щڣ(if��C΢Pi��T�/D�X�ӕLLj��a���3"�ِo-D�tiGl	�1f(�(S�t2��7D��A�L�u$�l�W��a�b�qm(D��2T��d�4U�WjA�}.�0��*D�@�,�~X6"�d�;;\H���3D���fk]Q�	��n_�x> p�/3D�$�sn��vL%�Q�I�s�r)T�/D�H�*�C��8ڷ���p����?D�Hsѩ��Dq�� �`��Z�"D���ԢC����B��1P4��?D���`��C�4M1�jK7y��9Pg�;D�\k�.��t���!�V]�~��g�7D�@�7m݉���6B� F0J�b6D� ˶&JEa�pQ&��_�.����4D����
0�|���ឞ}{���o?D���&�N'ʈ���l�@���>D�SS����#ٕb�B�H�>D���q�0(W�P�-Z�U��/(D��
&jџ+�u�)�.;���6`'D�K�������#��(�bL D����+K^T��M�&*��A�g"D� ��?=�*\1'D�z%���m5D�4��>->^�p�E�4Sq�c*4D����2Vlf�)2����W�2D��BE��NW���@쁓I���C�-D�\��&γ$�V�ږ�y#���+D��`��<s�������n��m3�Of�Y�$qJ�˄���$d�b�������M	F}��/A]Z=Psc/D��*�W5	B�hg��Z �b9D������Fڔ���A�,?M�]��6D�����_4c���kF�)�vŹA�2D��x���"b� Kp���,�he#�!2D��a���K��y���í�xY;P�/D���vC��&g��s�!�5G~V�k�;D���T��6���� �s�*U���<D���@��� �`a�!��J�q�S�:D��3JG�d'<�ME}� �
�h8D�����Y��=��HQ�`2���6�7D�T��[�
zɒ�7s��Y�$5D�h[�aǿD�@J�O²(�<���6D�{R���p{nT	�& ����@6D��q���ʆ���]�� mr�"1D�D�c^�$ajٹ�Z /~:[!:D��ZBl�	���A��2�V�P�5D�b�j�5���� �ɐZ0&l16�3D�ܚ�)vD�Q1��<Od���G,D�l�C˖0i��X�{�Rt�S�7D����)Rܼ4bR��K^�+G�8D��  A�$�#�l�Z�f ,��x
"O ��ِIRp�hM�M1�(��'3�����=M�Դ��c@��9�'���K����]��<p) E�'t��Х~��R#��>8��a�'��Mڷ&�N��ؑ��uBx��'�<{�%A�iu�Q��P�l����'��s�%��8��]����k^T�
�'�.U� �p̙�Dd�=c:i
�'����S�\f�$@b���'7�m�u��:Ut�)��G�g�Е�'^������=R��X*�$���'W*�[�ǃ%C+�����5��K�'M�`Ѓ9'2��y�n�&�R�'�����PZ�E&F"j`�!!
�'22�"�m��P���$_�|�	�'Z�$�P�P�p�$�KD�D3Gк-��'����Ҏ �-�|d"93J�)�'@N���@O%F8H#��+%@de�'�Y��Y�<�й��kL U��B.Y��C�#K{����bG�T�ȓ6;ڜ'�`�ȤO�#@��І�U��jg,�A�d�%a�w�8��ȓ&���5�ѻ�|�t�ϹAژ��ȓ�:)�f㖁'F< q2��ko����S)�U��d��u5fxJC�X X�4C�	3T)���"'˂R�`���	�2��B�	�	�m(�ȑZ0|Y�G�i�4B�	�X�RE���AP(�|W2B�	u*�
�U5�l����=B�Ɍ"ɰ�A�*_�q0���T��C�	�N���1���7��1���)��B�=C1�i���.�H��rdԶ�B䉖p�=`��gG�T{#�֔xJ�C䉈v0�$`�$Yc�D�a,��2�B䉿JӠ�І
KrL�4A��v�zB�I�`/�b�E�*:fV��?��{�"O��P�ަ����GBP01�F���"OR����(X6L����vo��X7"O�=�WM����S���qg-�"O~��BP;'.�M�F�%yOJ�g"OB��t����=���*=(�f"O��T�I��h��5
�ġ��"O4Q�V�]�z~����ڭn��z5"O��̶��(g͜�W���� "O�!���%l
�5(�Aȏh� !!g"O~XzB��' ���C�'��� "OY�,�J��ЂV�ŜR�<e��"Oԩ
���}/&�qB`�/Zy�W"OFdj3	�g%  .L/S$�dɀ"OP�2�D�yiHzӯʫ'��c�"Ot�'(
)h��2ϐ9
� ��"O��:��³u�z6�ڐz���"O��!�A�4�T�
��y���3"O�0a��� 9��I:��Ǫ[� q"O��׌��V7�3AjǸ�����"On�f�[8?�⁫�D3PY>�`"O��I#�AiR��*�&~hf��"Ov�)�-��Xd#dS6SM
]("OT5	0�X�v(�D��.K7^��"O,9B�"��L�H�m�\3|	��"O�p���W�kax ��ο?3���e"O��K�e��1B�����;+�ta"O���2�	9F�
�;�h��\��0y""O� B�R�
܁l�P�ٶƇ�H�ށhg"Oh��W$9�}
�Bo�BT�"O�P�@(4�>\����%{4�5X�"O��`CD_:e���tGԞR,�ju"O�@�'�=թPGI�$qk�"O����-]�R�8�F a�I �"O6y1f�I
A+2���N�J@'"O�!�%Cm00cE>G�4��"O�%ZB�¬mqz,: �Sm2�'"OL��e�Z
C� 9���J��v�s�"Ol�����^��0�hZ�}�.�z�"O�U
����4PҨ�	]��� t"O��4G�U�\ s.���tsE"Or��d��2��MU�n�����"O����DҶ,'�Y�'��QE����"O��#"�PnZ���Bڇ,�,X�"O2 �2�ܚ�:H�����4~!Z�"Oh�ʔD�
�Fp�T�8��"O�vϝ� @��U�0u,��t"ORV�U�` g&�����"O�ŐCI��4ґ�
8q����"O��@MɁ���(�bɴb�j���"OV��֠�zWl��C��!,:�$�""O�$��m�kH��g��	+(���"OҨk1i��j��d$�Q&tY8T"OL�qv�D�W�:���!2 �"O&��ŤF*Y�l�2������"O��Q�q-��3�mB��d�"OZ�r�� �
Dn�5x>^1�"O��2�L�F���r��10H�)W"O��4���T�N��E�߈/9<�R�"O�)i4aA�+���@���-��;�"O� �F.�:E6�̘�b��  ��a"O�`�����P�8u`OA�T*�)�"O�iD�Q�w8�ʡ�C�L�b��"Of�W�^:6"z�3@�6P���k�"O���� �2�X`��.���"O��!r�N�l)h$�?m#�qY4"O^���ɀ:n�`��''�,#�p��"O`	�"��9ڄYA�аVV���R"O�,QC޶X�`YSu�ã]Z�ū�"O�ݒ㢀�<>:�����yK���"O��ч^����s�ػPFl��u"O`q�$�L"����/40HR�"O������>ى���&,��"O���dіd��u��K���2"O�"�B� TP���s��y��X�"O }���']>�bE��g���[�"O&|����p��}�s#H�dy��9"O�Q��I�azh�W�I�yxn�H�"O�-HҠ.2�IЗ�P�1U�eї"O�ٸUg�38D<daPA\���"O ���3L�(��X!|���;u"O��ӗa(�����3pT���1"O��rE���z����A�ieԌy&"O�����ϫz�8�#�O[ Z��R"O
�;W�$�5+5/O�"I��"O8k���4(7�ذiZR�0�"O��"�͓!SSB��E+�<%:��"O> ��A�B�ld*E���͚c"O.Ɋ�����I�G�@5(:��"O�#��*�
 �P&؞t#^���"O\x�t���{��V	5~*���"OR��ß)6�8�qs�ZMd�Ч"O� ̥R)T�Ĩ��H� Z�BQ"O�H�&��`$�b2���Rf�02"O�=�B�`�����`D�,Lx��"O��k� ��ȱ�O�h����u"O��pa`O0/�>�+EoV�iۀ �"Of�d�j�en�x��,�"O�SS�΃[j�Z$@�!4�V�b�"O���B�)Xp�wN3 � e"O����h�=�ڵ`3-�;� �ir"OLԸ �"�|=g���=��U"�"O�y�c	���r�OX-<yj��t"O�Z"$EI�X1q�C�,V���"OkV~M��L�1Umj��u"O��q7E��s[j@�0D�/^b��"Oz�r5L�aZ�ax��^2�6Q�t"O:ĠLO�����#�(�K�"O�P֍��[��|�@�P1���J�"Oڱ�1K��b�
�N@�VT��C5"O�rDX�rX�����^6XB�"O��K�m�_�
�P�mM)7�츂"O�I��.���$ ЌW�~, �� "On�Id��u�\��K�:F,L��""ON�c��O�9ZH��)Y:C~"ܪ�"Oз�J�OĪ��y,"O��6��.t|�yQiE�?�t="O�5�4-�~��əg�Qm~X��"O�!{�h�C��Um��LTn�q3"O�u�r�� �VX5Nۦn7�8"O���ޢإSE$d ����"O6@yƩA�?�����P�%�:�r�"O��#�m�X��,1%A^�Na�"O�л���N�n	�c�0a`���"Oj�"��&}Nʨ9����c�64g"O��ug�\�9��Ƞ<�L�"O�a� ϟC�.���٩K�д��"O��PǗ)V���膱9id0"�"O�8Ȥd�(�`"��
�B{��b#"O���a�	!Y��s&FGPn�ق"O5Ʌ�Q<?m�9r�OH��0�"Op�Yt�=`�,�D�s��X�Q"Op�1/�<��c���2�a�"O�h{��
V�HT�`�41�1�"OE�]/6�G���S�"OV; n��k7h9�u/��4СX�"OFI�%O��HӺ 0�B�a�X�"O�W�A�ƭg�֐��"O�$�G�ī7�L��0�
���X�"O�f	�OL��ʒHF�JPN�
�"OP���Q�+�Z���gO�.*�83�"O ���_6,��ǲt��e"OĠ� �O*K�fX1^d4�S"O @�7mЯ�Dl�eĞ>����7"O a�Uf �dq>�O3�� �@"OQB+��s�b�{a�P���W!��= ��YibL�O�����K��VQ!�D�K���rf*R%Q<�KU��<l�!�Tj�MJ� ����JT�ŧ�!��^F�`�b놃d>6=i,K(�!�ą�dZ���^\<�y���V�:�!�W0U0R���,7Q#���⇣N�!�I!5�T�e(!<��� }:!�j5:�"'_ r����ǁX�9!�$
=f�,h�b�?k�DhJ㢞i!�dǹ��dxUD������ʻQ!�� 2]�q�I�969��l��P#28r�"O���G�h�@�5��Ό�uB%D���t�S�f���q�]����j$D�,�NG04����jW/Bɐ(�A�"D�4�t��9�fp3����^EP ��+"D�hHc�U5_d�;"��?]:�0�?D��9�ӵyJ�c��@%"�°&?D���Ե%�<}$k��,�0�a��*D���Ab�X枱��!ш0���'D��ʖȅ������O0u¬�Y�;D�����(P z4#�"4|�~���A9D�� ���=?�!� E
>+NzI�C�5D��Q�k��d����(
4(	�k�g4D���J��&�0�r�b ��as(D�hؠG�F@�0��A� ��Ae%D�,b��B�D!0 
 k2�@e�0D�$a ��0Ƃ ����!��$��g;D�(��6[�z��W'F�z>B�H&":D�x�IԬ���Ҧ�1v�C��9D�̘��m��D�Nޮ@��8D�ૅd�:�b�䯀�n5���׌6D���,W�|�X�k��B�V���2ů4D���voU�-i��AD��&~�\�A�&D�D�T��9m�}��G
F�� D� 0(Fm�� ƨW�d�(� 1D�(����E��@1c�I�x�8�)9D��K2m2n"]�"�u�@	8�8D��Fォdt�$�+���K%�8D����!��v���/��x�t
5D��Q�.B�%�(�r҆ %'�!�D��dAF�P�l�����rgf�Jm!�$N�T����l�$2Z�;�J�=GF!�$�F'x@�4A��a�b�"�I��$!��	2��=@v�� 48�hI:�!��ט2��"�#�Ni敺CȌ��!��ߥ��ՠ�+N�|YF���P�!�$�*S�0P32��pa$,�#n��u�!�ěa��B��y��P�U!k4!�ċ%�>����90�1���-!��Hx$5�`�c>!�$W�f�|0��׮���e��	(!�d�4q(�A�uB��(�P���"j!���?l�I:�Z�,�0��H�!�DH<p9�\j�����&@ϳ`!�DJ8��Y-1c��ӍI�u|a�'b���a�2LX��d�j�
1 �'̀�����S���83I��_Ǻ�`
�'ն�q�����)��g�^Q�q��'}���C�C�`�$hDA�C����'���рN��7t����=Z���'�*�S(�$Na�Æè�j���'\���#M>r�񃳢�39 P;�'�v�{_P���s$@W#`�x��'H��i��3��X�#���&$��'�:�rp/G�dLX�sc����a1�'Uࠁw�h��"���l��'���{ƣÂ�\�2l�=��E��'�㥭O\b�B.�R=��'/�C����h� "B' �0�'���oD;`��9��
�'I~隕Aҙ[X���A�נE>niS
�'
����8���[a�����	�'����F�7�JD�3mė}/h�(�'�Fi�q�D�� �E,	)������ ځ�/ґAt�s�c�Wz�۔"O�b�E@'@�pr5b��ʖ���"O>�wI��\����@��OS"]��"O~��#b��6]�0�H��,�x�� "O9X@f�1��p��&[0D�0����4S���$j���'���X?�r$ŋ�?ӂ��J�Q�6M!`��.=O�8q���?��
Ą`�0"�7��, .�V�6��.k>�P���3A�h�SH��
�X�m%�OB���a�ԺA؄Q`"�s�<�UDH�7\����|?�Aqf��d������'!R� ���?��d�ic.�TLD9���W��h�0F�O��O����O�p��늑8E*��5`�8V�P(A��'�7��O<6����b�� o�'�t���Iı'N�9�I9V]��0ڴ�?����?��'gS��p��?q�4��PID�!e����j��a 蘩5����(1�$��Q	<�֥�'�����X>μI�t�ӌ >
Q�'	�)e�7��/Q�P雐f9�"$QgcA�FoB��;�u�F)���ḧc���>&q)�!P8H,�@�iuH�����?9�O�T�sӆe�O� �؝��E�(4p��O��%�O~� ��8H�$U��h�K��<SW헱osfb����4�?��t�i�~�S��/b���G��:j@1�O����>
�+�C�O>���O0�$�������M3�(+��i�j@	{ ���lG�g��A����� a��ނK���0��O�� Dx���6p¼YD��8դ���h�y�ڸ.ua���MÅz�r�s�b�a��B}��6�TS�$��~a��C���f�c�؃7,��3V|���ȟDyI<�-���g��;�T�I6R��A[,��0�)�矠��NL6� Z��R�p�1�P���r�ҒO�ퟶʓc����2N�jI`l��� ��8@U���*a*� ��?���?	�G͍�?q���?I��:�M���YN�8V�.fp!�f��#������X ��I���Y�'A�}��f��~�P	n��Ȃf�6I�9S�*Vw�yu-��<z7�e��}�?i��Y���l�G�J%h�ꐤU$y��dx0!zǽil2Z��ã	�s�ӺӜO�v]�� �8����Ċr|�5Q	�'�>%B'N���e;`*�6c<L���'�66m����'�J���hb�H�D�O2�'#@x�K���V�(3F���X�0B+T5	��'�b ��ؚ�H�Ɛn|��Oқbnj��'+�t��ٝ3o\��_�a�d Dz'�	Vl���V

vp��۰@]�֝�N\d՛ i^�W��[�L0�$���[`��&������N|��4�5 �E_�3���j��ML���'L�O?��� g��� �ѕ.�ZI�#aE�@иD{���nj��'$��ݢ�+�*w�E ���J����?��3GX� ��r�t!��3(�'���n��`Y�,�������`����V�4��C�+�tZqK�,Ay�@h�I^����P>=���CIX�+b��lĵ���3�����@�A�H��Ɵ"Or�%	�%_��u׾�N]%?�ضe�D�3ͅ�s�=T��<�<7m׈yu��'>�6�O�#~nڈ+���E�&(
�er��c���I� �?��d{"ꁻ�)�?��(��jK%�Q����4�6��`���H�?b�"�r�ʣ~�M��#׾���=	�eT   �   ]   Ĵ���	��Z�Zv)Ċ;R��(3��H�ݴ���qe�H~-�8L,<���i�n�?
.Q�0�đmz(�Ӥ�._6��)�4<�>��' ��0O��@6�ʖ���:"m�&To�pS�Y2j��RߴZBqOR����D^*�MW�[	A�Ʃ+oY�Y��,���V���D 8Qf}I�4$���.�응e�:ל�;R}��c��e�Hu�Ҏ��K$ ����6)<��'���v�Z&(%�OR�2d��v�4�
��ȜJ���ʡ��g��o�$�?i�'Ed���=Q�)-O,��U'J�D��\c�(y�S菳tT,hĭG�WĂ)�O>��M8�zrF�O�mےl�&�,a�fg� M-BA<O��������OH�h2CS"g(�\�-�A��$�r�p�'��IExbkN}�)�?-|���!�T'.��Q�L���W��3F�D� )�����%ߖSjՙ��ʈ.
��J�A�'|ZuDxR���3�|PS�C�����tf6yӨm�}rBK�'�N4䧭<�rME�{�X`�b�,v~�l(O��9��D�<��'}l8�Q�20*i���5g� \A"�V~�'�%Ex��Vߟ�	wA̙D���1!.��8n��X!.&�I�8��x��x����w4����4zxӤ�\.�~R��x�'��(Eyr.ԱtCDI�s�M'�`R���?i$�d}B�8����t��u7:���*eB��t� GOR(�P�H�ƇN�7D,�O�%���\�'}����C]~��t#��� g͌�	4��M>�d�ۈ*6�Q�<�I�)�Xa�(Y�=lT�fЯ�PX��'Nl��@ ��"O��Y�N-W*`���R	Hܩ�D"O��h�f�;P�&�@2�"x�a�3O��x��� K�JQ���ʤl������f���D�4�O�jR'�j�V(�l�P�.��u�	�]�9r��B�T��O:���b�F�44X�(v U����'Q�����3!pĸ��EY�N��I��O��C&��,��l�m
T>��¦��@t�r�lF>]���pH5D��"�/[(j��	���Ĳ���YRL�/O،hVc��9:`<%>c��;��&���į�%!Fb1�-'�O���פ��]i�]k�f�:�%KPN"�í2���B�'�~}i!`�'j[+��I&A�����)��X�KY[���O�q)T�ڱD�� s-�E��-��'aL��⊯\�-3%�>�fix�Ox�Ұ�X�/��If�[>a�    �    R  �  �  &&  x'   Ĵ���	����Z�/C�'ll\�0�|r�'a�	�Dط8��0b�
�<�}#�'�t4��B�h�dt,�:?������i"x�	�-��K����1Bʚ�HH�� Ҕz�J�[�.�0�|)`��u䨉:�Œ�_2Ii�$]�-��s�	��	-�i�V���LX��92��6�x)����sA�)(E&X�9צ��
����q�`˯do���ЂL99}�4y2�E�C����>��(J�"���U�i�����m�<�e���Vk�$�r���3�,���E^�<�Ѝ3?�0���x"���,�]�<�BcQ�P�nЈ�"R�	cT����M�<YDc�r��1��Y�����F�<Q�ձP�҅����*
8�P{6�B�<鲆
(z8���J�%~A�C�N_�<1�!+��|�p!O!gƖkB�F�<��o	�;��B��[;Q�xYq��~�<�և�+}xe薋���b��d�Qf�<�!��.0� �a�=5l���
d�<��"Ι%yMX$(��^W$���|�<I$l[?E~*�l�!Ha�T�C�y4xF~8i�bL�qȂp���y�)�	{O�|���
�txf���J�ym �}Y�*#*��7\�@V$C7�y�M+,:Ѐ�JB�9�0C�gN�y(�q�:�$�M⧄VG!�T'!w���3�X,B���]!�LJ�.h�wD	�6�a�P��(v(!�D4 ���H�o"ʁY��ѻt�!�$!W[V��1΀! 1��F_Z�!��T�Ms�@�/��j���wFòk�!��D��(��&o��B�/E�!��q�%��O�2�&yz�΅�k�!�D��6��<	o�R�(�`�M�<!�ĜRq���Wc&V��K�-<!��yy�����b$�Њ�t/!��H�fؠ���0�����V9!�C�p}܈r�j��Se<���Α�B䉭W����KD��	 �3|pC�"Oh�q[�	 �j�h]j5�փO-�C�I�"�� �S������0��C䉴([4��BH
C��]�2���1˨C�I�3��c0�N�j��q��&����C�ɸ���[2��1-�Q&�̧:�bB�I.t*�]�7+W(8C�[�/Р"�2B�I�r�@�D ���H2���
B�UCL�⋀2:*�b�;|�C�IRU@��m�	8���k��M�BB�	/���ck�u���"D��!:�C�	8W%����o c~�E�D�î�C��
=�x�0�E��-"0�ˆ��7D�fB�	�+���ħ�bm�V�D�y�hB�I;=���+� >�@�1/�4+%XB�	�~0��ԧ�3[i.i�0(��sxB�I,\ ���d�ѵ3!b���S�BB��9�0H��� C'��Bh��)�C�I\���ao� �Ď���C�	;A�d5`���/}����C�(%�C�ɯmh|dZpe��o��0��-�eA�C�	��f����N�h�\�'F�B��C�ɣ;���{LG�s�r�
fσ�l(hB�I�v!��đ$8)F��� �Ju8B�ɣ�dX�g$�6%"��P�S�&Z�C�	��PE�e3}�]�g"ݯ~��C�I>�a��"�1zr6���"X3ZB�I!^0���"#�-<����DX�L�B䉛jwL��JݳM]�X%��`8nC�)� RL�6g\�F�
��f�%Z�"OmQ�2����w	I.80��"O����,���"��c�N�3"O�U��M�B��L�sȞ�M_r���"O��V�>n�A�l&X]+q"Ox In�>�j���	��v�lA@"O��Ct��C�����4E�f�+E"O��1�ED/Cb4�����`)1�"O(� ��bR�@��0���1"O��1BոL�|<"<H�Hq� "O�k��&S<EQ��-���%"O� AqВZ�RP�%����S�"O���cLa6���\Ȉc"OJ0� &Q�z��@I��[�_|��"O��V���:C�t��GB�U�p�i�"Oͨ�k�7���s'��1�U[a"Ov�+v-N3�j@��e�[ߚl� "OZ�b/2�tC1�M�dȞE�r"O8��O�#3�)YE�R5`|�e"Op�ʖA���8�f	�}���"OB�xT�L�P�a��7�%!�"O�8ش��)��t��닦,c�}�3"O�)��M͜�� ��JկZ]�3"O(���	�*�\XtI�xJx��s"O�Y[&�K�AT%���E����"O�-��-Q0 ���K@Kۨ\{XS�"ON9�F�'Tࢯʿ;Q$��"O|Uc؋e$�r� � V��}��"OHp�)��.�a�
�%O�� "OH���DG
�B4�q�L?D�<�*�"OJ���
.q�u
�9�>�s"O�K�%\,NHw	ή8����"O6�˗�SfT����/
��h��"OR5�A,!L2��OS1s��3D"O>q�&I�D2��bNح)���%"O��F��1&ʄ�#��t�#q"OX�����IZP�����3�X��"O^�U��ZrΔ��D���"OL�auGH�|�P+�Ů���"O
���Z3R����鑘b%Ъ�"O���*��? �	�hcܬ��"O�{U�;ø$�ceH�e.���"O�)��ٵj�����Q3'V�@�6"O��Ң$B�O��X�j�ܑ�S"O�Ds���4��R�hN�C��D�G"O��U�O
.1���SD�2��"O�$�R�?OH$q6/ҹ~0H0��"O"�SGF\=RY�#�A&�;�"O,hRe��9Lv�]�%�������"O\�s�M�W��	1��)�BP:'"O
y��D��-$�S�0e��Xxc"O��"�'I�pZ~=2�N�:�6(�e"O�1�7Y�i�PO��85����"O�)��͂&�ikw͕9#�2	�r"O���@�R�������'�,�i�"O8ɱa�٣g��U(sA@�t��e��"O2��SƐ(/9�]ЕG��I� 4�"O ��5������&K�h��\�v"OdiD��"y:�3�>*�"O\�K1�H�]
���
:<�P �"O��X��3�f!CvkFq�d[�"OD������RA^��ֈ$�"O������B���sf�G䨚�"O���Q�Y�8�
�{`�϶X1��ڀ"O� <�G�S/N��0��3M�,�R"O�T%*��x�V!z���|��"O�$r�)��=�l�j���
0�2L�A"O8���I�hV��  ���0�.�c"OT9rn��.�{h��e����"Oe�&o�$t*8Y1�9b��"�"Ot���6���b���bVb�XG*Of���̌����h�H��m����'9:ٚ���-�T� ���P���'�hiC�����K�^0�	 �'�>�bH��^�։8`���R�v=��'��5C���t� �:�ڶi�'��@feC,Sf�P���6F� ԋ�'�t�jb凌0��=Yu��Ky��
�'�pB����<4�$	�,O�Y �'P��c�a�7u�,��ۋ
!F��'Z.@3拌5gf%xg/ܟ h1��'�}y�)Z�=$!r�E�A�4�p�'��xx��o�& ���(w���0	�'ђ]yA`�)"N��"���Z�Ν
�'Q�������!��O�_�* ��'����a&N�{���ѷBR�<�'�@�0�c��,#PQ�4,̋L�x=�'�(J ̊�.�@[�`��~X�`	�'�d=`2��R	�mkƃ��w�+�'��� 針ϊ��1�OOTC�'�6�pED[�.�bp�ƌ�X2]�
�'� Yi�%;
*��E�/_k���'�hu�Ǭ	!f��,��a�G��\�
�'Z�T��x���U��͉�'H��#����xИ$�U_	L� �'�z J�*�&j7�ˤ@�6W��;	�' 
u�E��& ����"Ҍ]	z-��'TDQ{�!��_ H��9b�8�'�Xbc	4qw����!�Ϩ��'� �CmK�o�`��g����A��'��)(Eg?z��-�!˻5��mQ�'�<��Gˋ�[�H`��З7'�t�	�'��Hr��33Z�J�a�>#���P
�'@|	H�i2yN�@b@��1�	
�'�B��e�{�vlx������'�a�v!�+�Is�̝�Y
�'��djG� }��Y��K��3�'�v)�!i� 0��́r��$t��	�'L2���B��(�`'� � �"�'ir@�*M<nh��+Q��F` �'�nL�A')���ĉH?����'�d�`�"˘?+�� �h��<���
�'��q0��Ǣ\f���7���3Ϭ`�
�'�f�[���(U��`����#�$[
�'(̪�E�.\ԡ�1
L���j�'~E�s(*�ԋ���O�f���'��yp N�%f�ơ8$�ͧo�`"�'�49�i_���E䋘�8)����']�u{�l� �*�ɠ�3>1��'c4 v��@�T�JC�:�X�B�'� ��K�/��)�s�*9�\�	�'�$�
E`��1�tAYC��(t�	�'�0�j�D#H�<�ӌ/)��tY	�'4�C,O�=�<�g+׊5/���'4)ˁ��,։H��5�`���'X�4���X
G���iB*�o����'>��r�֊.���u����5!�'�A�(ON����NJˤ�+��� ��H��"4	�	۸rb��t"O9iE^�U<Mp֯ϲ=��� `"O�\�v ��0��E�3��\�"80�"OVI�
[�8p6MYG*�<X���"O�a#�+�o�H���F��Q"O+M��l4́1fO��{��W��!���:B���H�"A�ls��ޮ�!��T��*1�	D(y�(e�!���7 ������ß"c(���ʝ�;�L|�Z�����	�U���A0f��M���z�AS5}߈C�ɨ_��y��$��諤�;GO�B�I`�l�s@�"i��C��B�Ɉc]NL	�Y<,p>��B͍!_ B�I�"(����;�J�*ׯʈt��C�I�'q0҇KL�k�Dl�%���7%�C�ɘa6x(f-T��!I�R�JTB�	�no����N<J_ar�D��$)�C�I�~��D��A�$9X�H�3:�(C䉛62l�����:Qs���2A]t8C��
�QČ�uH�m�����4C�ɰ4,�9��/�}�DS��8HC�I:s*�$sB��}��M��	۬<XB��	) l�
�ϗ <TԽʁ�ܝ�\C�ɰw�,02��"M�dq-�#qC�I%A�4��2��=���a��U�[l2C�	kS�"ң?D�9�%�&V�C��#W�
e�aS=)R`�	`�`,(C��
����c�@9H7�1��+�L��B�	�7�V4��KD%���₢͇*��B��pT\���7bJIR5Ν,U��B�ɃG��8�3�WvP�ȳǫ�u�ZC��C�va�pIW6IfX�Y��G���B�ɯ�
���N�:J2&Ѐo�r\�B�I�Y�d����<#d��$�8D�\C䉾7ܴLRG�§:MrӧN�q)^C�I�>e �b,ؘld���a9U�B�I1>�,��<��T�eFL��~B�	��ؘd��l����i˅�xB�ɯwc``BƊ�9j�p�� ��>��C�2do�X�B���d4�u�˙nK*B��#Q��E�E�V�A)<*��\�g�(B䉁R��� iؿ6�+fě4B�B�$\�� ���҃B����M3�C�	L�f�2v!˙{+*����6{&�C��'^������U>Č:a�ȵ{
�C�ɹy`Jpɒ��	d׆��0��2x�C�2w@v�CƬ�-�\�+�f��D��C�0b��a��ϑ4���`�	y/�C��h��b�A9`���;ׂ_&"�LB�ɖ`���p��^33<xu㥍><�&B�	��Eb�J.z�H��h	�y��C�)2�H��L�Go�Q��JC
M�C��<C����E��N ���l��C�	�\<N��#�G�9�n�!���[��C��2w@L\9p'�!&n:�t@�t�C�ɸ�0���H� �5�h ��"O�1i��$a1�%��N#���w"O��။�=�;�N�dnI��"O4��1cM�{jY;��@�~4�[�"O����+U2�>Ds�,1�(�D"O�,��d,
� �LU�e�h��"Or�X7��'�Th�����Ф�e"O��
��ݫ*|�!�*_�{p��"OV���mځ-(Ah���fĭ9�"O� ��Au��!pe�r�#VmC�m�"O��B&D��qQd#)�졐P"O>�&���T�
	�b^t��E	�"O�������l��YG�&���"Ovѓ1IZ�~�B���<���"Or\�Ԉ��Q8��Ǌ!;�"�Ѓ"OL��"A��^�|���}�̴��"O�(��*ٵ5Ȳ]���="1�5"O���#Ip�Q2��E�1�"O�Yk�d��CtCƣ�tzd"O�B���:�d��vǏ��~�"O^�h��!�0�r�EQA�|ZT"O�e�b�Z�E�X�7ś�0�v�;�"O���קÇ ���c4��3	nd�H2"OA���D:]�:�+�dC�WevВ�"O��鐀љS�&�1vAD�j>pd�w"O�Ѱ7O����V�X#���%"O�|�$j�{[`��$��K�80�'"O��c4&ǆuw��'B� j����"ON=�/B�H�ോb� M�1[g"Or�
e���ޕzf���5�
ŨT"O���g ���}�a��6���[�"OB�Z>]����ɋo&lA5"O��2�.ɥ"��E�'��8&�H"O
�O�!|1�$���5W�8S�"O���皅t��p!	K�����"O�(���L}����+D��}h�"Oj`"��
�4YR�VO�"J��"OF]�f'J�~{���Q��-j��"O �#$jJ�& �1t,D�o_��(�"O�$��Z� �:�+��$<:�S"O��Z��7"M �2�X����"O�0rfhR;j��T FfE,�� pt"O<Ձq�٣<a��Җe��|��)8�"O�Q`i��~�˳N�M��E��"O�X��]!j�z�ʲg�$���"O�RQ���:x@�&旯Mΐ�%"Oh83���u���@��1r�b�+�"OBU�&e	�Wr�c5��rߊ%�d"O�[V%�	�00���NΞQ�"O�Ѳ3o[a�D��?mZ�*f"O$�V��/?j�A5BO�gNr�a�"O�Uk�e�xz��O�6C�I#�"O�����״��狊�ba)�q"O�����r8�r��5X����"O����Ώ�*dX�RIƀ@T��`1"O@R�+cq~Sw�֨_>�i�"O�ɘ D	T@��� ̯Tŀ�		�'�J8�Fo_;iQ��HS
�b9�'A*���+�
Z*�S� ��>�+�'�:�u�
~j���rg��	ޤ�'�"�b��$KU,t@��M3���'��8�H��dK��Q1�^~
@��'�hh��Ȃ���yc�ȶ�nL��'�(���8�ԅkU��x���K�'�P8��
LAk���.��h��`!�'��j��^+q����dgN^�4�8�'`�A���{��e񠝉P��h�'=b����b��%
Q�]�LRFD��'���Z&�@G(TK���G� �
�'�|�����<�8� #�P�r���'���5� [�p�oQ
	?Ҩ��'��iD�������E��t��'���hAe�0{A�]�@!��s�"O� ��it�̮w�X#��U�i���p'"O<���F]�h�H����E�)�
#�"O�H2�� &�~ŃW%I�i��8��"Oּ�Q~AZ��A]��M{�"O2`����;�e���<?v&��"Oq@
,0�H���9���r#"Op���h�R��%͜A�X�4"O�bdm��.�n :��¥w|N	sa"Oȅ����~8ȡA1��q�A��"O��S�R�@Ъ�����! X��I�"O�u� �0f�Z=�ꗆe�
pb"O���G&ɶc;���J��t��<��"O�Q�ggd\��(ң=�zm�"OL1���>V���Є�D�bΦpa"O�lS�m��?����W�`�
��"OPy��7	r,P���"�xʆ"O`�������X�=��Y��"OT�ڥ"�*\xi�� g{�,+c"OP�Pq�C�F.6�Z'��^���i'"O�����<O��Ex&�Z�Cy(U˅"O������z��鳒�!<O`�Q"ON���O'Fp����Ȥ[6�-XP"OJ0ˁb�>(��ظE)��T��U��"O�Ȁ�+��*�*%ZI��w���R"O�	
���R��D������c�"O���!ڸ��q*�ǋ�`����"O�䂐�@z�܌���K#����"O0��"��(Ј�j0-º� T"Obh�r�.+�0C����,E�̹q"O�S���|ء�&�$=�}X "O��R�?��[a`��/:� �"O<�;� �=��4�q�_�&��"O�XǤT�t�\A9E�ǒy�혰"O���N� /�0IA%G�u�Yv"O*c�&�t���r�B�T	� �"Oe��!�$9t��f�_�"�|���"OR`rv#LHH�I�i�4B�pLQu"Oڽ���� ^��E	�~�p��"O��AG
�>�>d��g��� �"OB����[�P��d� fU �=�"ONI,,��"Q�**a�*[�!�d�7:�d�V�Q�~�6����T�D�!�Z�A�ܵ��m�	E�bO��!�d��l2��#+�2 :�`��� �!���46(���J&P�y����	W�!��P�o�vMZ�B�|��1���!�C>^�X���{��=��얖o�!�ă�<ۼ�2f���I0=�JD�e!���(A�^� 2�Z�F�l�K��A��!��;wA�\�ש,H�� b�@5!�ϓ(����m�09�P`˽q!�D@�Gl���]�O��`g�1m�!���r5a%+°L{��1�Ơz�!�D
�;@X���N,�[���Q!�$O��$����b�ڠGX�,a!�f� ��X�~_�mA&@�$!�D���l5�#�JW���q���>!��/zV��I��mSԂլ��u!��^�rh����=q��sDMZ�Z�!��5Rz"@�����6DJ�Z
&�!�Ԅ8j  �d'�4D���F�!�$];��!4M�p���Sc�V$G�!����5A&O�R)>=q0$�!�d�6tF�cB�;r�Yc��j!�� �$c D�u�ʌ@�R�5/f�s"ObP�����C"��:P���*�0�`�"O�9�J��:�H�;��&U�
5�P"O���^XI�����9��"O��X&�֕F]�Dm��`=�"O�ŲEK�6=a~ɲ���!J�{�"O4\ɒ��-+V!��%g�#"O�%c�Òr di�Hج<|��"O�� �鄌uܘ�'��O�|�"O�t�/�R<p8���9�@��"O��QV�D�*>�h���"����"O�|Cq
�1�t��$i	(P�zM�2"O��Ы��)�q�Gǉ�SbF��"OB���  �   j   Ĵ���	��Z�RV)Ǒ7>��(3��H��R�
O�ظ2a$?����H�49a��i��I��i� ]�=����V`�6̀��9X�4Z���a�'[�V��p�4�I�8QP�Z�d��V}@����2Sd#<G�5x�67�]�|mN![g
��{� < gÌ,%���`8����2��L�OUrQ��_�qJ��'h�As&N���3�f�p4�+��5��L�?{�L%�z#
1;w�Z�.���ԟ6��6D�	2K�*ְ���qn<!(��C�+R!" �O�� �%�W`6�h�X�����<���� D�>b x�֍_�Ԓ�-[�2$R��'׮���d	@�'���'�)��N�6"� mԈv,�4rhe��i��I"5��H�/X)c7�!B-�2N$K' 8�O���Ď#��� [��e�@X1$s�����L)tg�H#<��6�Iƒ�l�D�<\:��iМ�B��i�qDx�k�L�'�t�dW5@eĸ3ڳ<=��IY��'pz�Ex�p~�JÝi!��p�A�Q4��[5�ի��$�'�O������,-d�FB��L�2�H��خ7�4Ex���f�'D�!�I#e����0fZ ���C�6h$�b�( G�I�'{0�PrNЀv�(0pC�D�441�'}HDx���I8[���fKG?�d��fc��e���T�ۚ,>� �%o��Y+ߴRk�|CCJG�'t��*����u��ߢ&XTx�@�ڈI�DX۔
�^qORl���[
����X��ǈa� �:Ή�7�P��%X6�q'����(O<U��ҳf����Ϩ(2���"O,���  ��]�\	.#�p�A*��Ɇ4`�(�b�V����hR��LmJ��B�&��G=�¡:Wid�E�CF"t�p�җ#�3u�	���M��$@# �<��h
93Q�����-A"Kc�\�"�O��0«?D�0�k�%k�r��"T�]v�ʀL�<��'�B�0gTd
̀1႕19J"ܮj�FDB�'m���@��|ɠmҋV&X��דj�2i��)b��;����F�H��3?e{�N��2W��# b�Gٹ_�<A��cy���3�j��M(����$���	�� �=��$ ̐P��gR!:��I""�L|�#h�29�B䕴f�y��_�C:9��#���?Q�HA*1��J�\?��,p�e�����4����ݲ�(O�t��S��,
�8    �    R  �  �  &&  x'   Ĵ���	����Z�/C�'ll\�0�|r�'a�	�Dط8��0b�
�<�}#�'�t4��B�h�dt,�:?������i"x�	�-��K����1Bʚ�HH�� Ҕz�J�[�.�0�|)`��u䨉:�Œ�_2Ii�$]�-��s�	��	-�i�V���LX��92��6�x)����sA�)(E&X�9צ��
����q�`˯do���ЂL99}�4y2�E�C����>��(J�"���U�i�����m�<�e���Vk�$�r���3�,���E^�<�Ѝ3?�0���x"���,�]�<�BcQ�P�nЈ�"R�	cT����M�<YDc�r��1��Y�����F�<Q�ձP�҅����*
8�P{6�B�<鲆
(z8���J�%~A�C�N_�<1�!+��|�p!O!gƖkB�F�<��o	�;��B��[;Q�xYq��~�<�և�+}xe薋���b��d�Qf�<�!��.0� �a�=5l���
d�<��"Ι%yMX$(��^W$���|�<I$l[?E~*�l�!Ha�T�C�y4xF~8i�bL�qȂp���y�)�	{O�|���
�txf���J�ym �}Y�*#*��7\�@V$C7�y�M+,:Ѐ�JB�9�0C�gN�y(�q�:�$�M⧄VG!�T'!w���3�X,B���]!�LJ�.h�wD	�6�a�P��(v(!�D4 ���H�o"ʁY��ѻt�!�$!W[V��1΀! 1��F_Z�!��T�Ms�@�/��j���wFòk�!��D��(��&o��B�/E�!��q�%��O�2�&yz�΅�k�!�D��6��<	o�R�(�`�M�<!�ĜRq���Wc&V��K�-<!��yy�����b$�Њ�t/!��H�fؠ���0�����V9!�C�p}܈r�j��Se<���Α�B䉭W����KD��	 �3|pC�"Oh�q[�	 �j�h]j5�փO-�C�I�"�� �S������0��C䉴([4��BH
C��]�2���1˨C�I�3��c0�N�j��q��&����C�ɸ���[2��1-�Q&�̧:�bB�I.t*�]�7+W(8C�[�/Р"�2B�I�r�@�D ���H2���
B�UCL�⋀2:*�b�;|�C�IRU@��m�	8���k��M�BB�	/���ck�u���"D��!:�C�	8W%����o c~�E�D�î�C��
=�x�0�E��-"0�ˆ��7D�fB�	�+���ħ�bm�V�D�y�hB�I;=���+� >�@�1/�4+%XB�	�~0��ԧ�3[i.i�0(��sxB�I,\ ���d�ѵ3!b���S�BB��9�0H��� C'��Bh��)�C�I\���ao� �Ď���C�	;A�d5`���/}����C�(%�C�ɯmh|dZpe��o��0��-�eA�C�	��f����N�h�\�'F�B��C�ɣ;���{LG�s�r�
fσ�l(hB�I�v!��đ$8)F��� �Ju8B�ɣ�dX�g$�6%"��P�S�&Z�C�	��PE�e3}�]�g"ݯ~��C�I>�a��"�1zr6���"X3ZB�I!^0���"#�-<����DX�L�B䉛jwL��JݳM]�X%��`8nC�)� RL�6g\�F�
��f�%Z�"OmQ�2����w	I.80��"O����,���"��c�N�3"O�U��M�B��L�sȞ�M_r���"O��V�>n�A�l&X]+q"Ox In�>�j���	��v�lA@"O��Ct��C�����4E�f�+E"O��1�ED/Cb4�����`)1�"O(� ��bR�@��0���1"O��1BոL�|<"<H�Hq� "O�k��&S<EQ��-���%"O� AqВZ�RP�%����S�"O���cLa6���\Ȉc"OJ0� &Q�z��@I��[�_|��"O��V���:C�t��GB�U�p�i�"Oͨ�k�7���s'��1�U[a"Ov�+v-N3�j@��e�[ߚl� "OZ�b/2�tC1�M�dȞE�r"O8��O�#3�)YE�R5`|�e"Op�ʖA���8�f	�}���"OB�xT�L�P�a��7�%!�"O�8ش��)��t��닦,c�}�3"O�)��M͜�� ��JկZ]�3"O(���	�*�\XtI�xJx��s"O�Y[&�K�AT%���E����"O�-��-Q0 ���K@Kۨ\{XS�"ON9�F�'Tࢯʿ;Q$��"O|Uc؋e$�r� � V��}��"OHp�)��.�a�
�%O�� "OH���DG
�B4�q�L?D�<�*�"OJ���
.q�u
�9�>�s"O�K�%\,NHw	ή8����"O6�˗�SfT����/
��h��"OR5�A,!L2��OS1s��3D"O>q�&I�D2��bNح)���%"O��F��1&ʄ�#��t�#q"OX�����IZP�����3�X��"O^�U��ZrΔ��D���"OL�auGH�|�P+�Ů���"O
���Z3R����鑘b%Ъ�"O���*��? �	�hcܬ��"O�{U�;ø$�ceH�e.���"O�)��ٵj�����Q3'V�@�6"O��Ң$B�O��X�j�ܑ�S"O�Ds���4��R�hN�C��D�G"O��U�O
.1���SD�2��"O�$�R�?OH$q6/ҹ~0H0��"O"�SGF\=RY�#�A&�;�"O,hRe��9Lv�]�%�������"O\�s�M�W��	1��)�BP:'"O
y��D��-$�S�0e��Xxc"O��"�'I�pZ~=2�N�:�6(�e"O�1�7Y�i�PO��85����"O�)��͂&�ikw͕9#�2	�r"O���@�R�������'�,�i�"O8ɱa�٣g��U(sA@�t��e��"O2��SƐ(/9�]ЕG��I� 4�"O ��5������&K�h��\�v"OdiD��"y:�3�>*�"O\�K1�H�]
���
:<�P �"O��X��3�f!CvkFq�d[�"OD������RA^��ֈ$�"O������B���sf�G䨚�"O���Q�Y�8�
�{`�϶X1��ڀ"O� <�G�S/N��0��3M�,�R"O�T%*��x�V!z���|��"O�$r�)��=�l�j���
0�2L�A"O8���I�hV��  ���0�.�c"OT9rn��.�{h��e����"Oe�&o�$t*8Y1�9b��"�"Ot���6���b���bVb�XG*Of���̌����h�H��m����'9:ٚ���-�T� ���P���'�hiC�����K�^0�	 �'�>�bH��^�։8`���R�v=��'��5C���t� �:�ڶi�'��@feC,Sf�P���6F� ԋ�'�t�jb凌0��=Yu��Ky��
�'�pB����<4�$	�,O�Y �'P��c�a�7u�,��ۋ
!F��'Z.@3拌5gf%xg/ܟ h1��'�}y�)Z�=$!r�E�A�4�p�'��xx��o�& ���(w���0	�'ђ]yA`�)"N��"���Z�Ν
�'Q�������!��O�_�* ��'����a&N�{���ѷBR�<�'�@�0�c��,#PQ�4,̋L�x=�'�(J ̊�.�@[�`��~X�`	�'�d=`2��R	�mkƃ��w�+�'��� 針ϊ��1�OOTC�'�6�pED[�.�bp�ƌ�X2]�
�'� Yi�%;
*��E�/_k���'�hu�Ǭ	!f��,��a�G��\�
�'Z�T��x���U��͉�'H��#����xИ$�U_	L� �'�z J�*�&j7�ˤ@�6W��;	�' 
u�E��& ����"Ҍ]	z-��'TDQ{�!��_ H��9b�8�'�Xbc	4qw����!�Ϩ��'� �CmK�o�`��g����A��'��)(Eg?z��-�!˻5��mQ�'�<��Gˋ�[�H`��З7'�t�	�'��Hr��33Z�J�a�>#���P
�'@|	H�i2yN�@b@��1�	
�'�B��e�{�vlx������'�a�v!�+�Is�̝�Y
�'��djG� }��Y��K��3�'�v)�!i� 0��́r��$t��	�'L2���B��(�`'� � �"�'ir@�*M<nh��+Q��F` �'�nL�A')���ĉH?����'�d�`�"˘?+�� �h��<���
�'��q0��Ǣ\f���7���3Ϭ`�
�'�f�[���(U��`����#�$[
�'(̪�E�.\ԡ�1
L���j�'~E�s(*�ԋ���O�f���'��yp N�%f�ơ8$�ͧo�`"�'�49�i_���E䋘�8)����']�u{�l� �*�ɠ�3>1��'c4 v��@�T�JC�:�X�B�'� ��K�/��)�s�*9�\�	�'�$�
E`��1�tAYC��(t�	�'�0�j�D#H�<�ӌ/)��tY	�'4�C,O�=�<�g+׊5/���'4)ˁ��,։H��5�`���'X�4���X
G���iB*�o����'>��r�֊.���u����5!�'�A�(ON����NJˤ�+��� ��H��"4	�	۸rb��t"O9iE^�U<Mp֯ϲ=��� `"O�\�v ��0��E�3��\�"80�"OVI�
[�8p6MYG*�<X���"O�a#�+�o�H���F��Q"O+M��l4́1fO��{��W��!���:B���H�"A�ls��ޮ�!��T��*1�	D(y�(e�!���7 ������ß"c(���ʝ�;�L|�Z�����	�U���A0f��M���z�AS5}߈C�ɨ_��y��$��諤�;GO�B�I`�l�s@�"i��C��B�Ɉc]NL	�Y<,p>��B͍!_ B�I�"(����;�J�*ׯʈt��C�I�'q0҇KL�k�Dl�%���7%�C�ɘa6x(f-T��!I�R�JTB�	�no����N<J_ar�D��$)�C�I�~��D��A�$9X�H�3:�(C䉛62l�����:Qs���2A]t8C��
�QČ�uH�m�����4C�ɰ4,�9��/�}�DS��8HC�I:s*�$sB��}��M��	۬<XB��	) l�
�ϗ <TԽʁ�ܝ�\C�ɰw�,02��"M�dq-�#qC�I%A�4��2��=���a��U�[l2C�	kS�"ң?D�9�%�&V�C��#W�
e�aS=)R`�	`�`,(C��
����c�@9H7�1��+�L��B�	�7�V4��KD%���₢͇*��B��pT\���7bJIR5Ν,U��B�ɃG��8�3�WvP�ȳǫ�u�ZC��C�va�pIW6IfX�Y��G���B�ɯ�
���N�:J2&Ѐo�r\�B�I�Y�d����<#d��$�8D�\C䉾7ܴLRG�§:MrӧN�q)^C�I�>e �b,ؘld���a9U�B�I1>�,��<��T�eFL��~B�	��ؘd��l����i˅�xB�ɯwc``BƊ�9j�p�� ��>��C�2do�X�B���d4�u�˙nK*B��#Q��E�E�V�A)<*��\�g�(B䉁R��� iؿ6�+fě4B�B�$\�� ���҃B����M3�C�	L�f�2v!˙{+*����6{&�C��'^������U>Č:a�ȵ{
�C�ɹy`Jpɒ��	d׆��0��2x�C�2w@v�CƬ�-�\�+�f��D��C�0b��a��ϑ4���`�	y/�C��h��b�A9`���;ׂ_&"�LB�ɖ`���p��^33<xu㥍><�&B�	��Eb�J.z�H��h	�y��C�)2�H��L�Go�Q��JC
M�C��<C����E��N ���l��C�	�\<N��#�G�9�n�!���[��C��2w@L\9p'�!&n:�t@�t�C�ɸ�0���H� �5�h ��"O�1i��$a1�%��N#���w"O��။�=�;�N�dnI��"O4��1cM�{jY;��@�~4�[�"O����+U2�>Ds�,1�(�D"O�,��d,
� �LU�e�h��"Or�X7��'�Th�����Ф�e"O��
��ݫ*|�!�*_�{p��"OV���mځ-(Ah���fĭ9�"O� ��Au��!pe�r�#VmC�m�"O��B&D��qQd#)�졐P"O>�&���T�
	�b^t��E	�"O�������l��YG�&���"Ovѓ1IZ�~�B���<���"Or\�Ԉ��Q8��Ǌ!;�"�Ѓ"OL��"A��^�|���}�̴��"O�(��*ٵ5Ȳ]���="1�5"O���#Ip�Q2��E�1�"O�Yk�d��CtCƣ�tzd"O�B���:�d��vǏ��~�"O^�h��!�0�r�EQA�|ZT"O�e�b�Z�E�X�7ś�0�v�;�"O���קÇ ���c4��3	nd�H2"OA���D:]�:�+�dC�WevВ�"O��鐀љS�&�1vAD�j>pd�w"O�Ѱ7O����V�X#���%"O�|�$j�{[`��$��K�80�'"O��c4&ǆuw��'B� j����"ON=�/B�H�ോb� M�1[g"Or�
e���ޕzf���5�
ŨT"O���g ���}�a��6���[�"OB�Z>]����ɋo&lA5"O��2�.ɥ"��E�'��8&�H"O
�O�!|1�$���5W�8S�"O���皅t��p!	K�����"O�(���L}����+D��}h�"Oj`"��
�4YR�VO�"J��"OF]�f'J�~{���Q��-j��"O �#$jJ�& �1t,D�o_��(�"O�$��Z� �:�+��$<:�S"O��Z��7"M �2�X����"O�0rfhR;j��T FfE,�� pt"O<Ձq�٣<a��Җe��|��)8�"O�Q`i��~�˳N�M��E��"O�X��]!j�z�ʲg�$���"O�RQ���:x@�&旯Mΐ�%"Oh83���u���@��1r�b�+�"OBU�&e	�Wr�c5��rߊ%�d"O�[V%�	�00���NΞQ�"O�Ѳ3o[a�D��?mZ�*f"O$�V��/?j�A5BO�gNr�a�"O�Uk�e�xz��O�6C�I#�"O�����״��狊�ba)�q"O�����r8�r��5X����"O����Ώ�*dX�RIƀ@T��`1"O@R�+cq~Sw�֨_>�i�"O�ɘ D	T@��� ̯Tŀ�		�'�J8�Fo_;iQ��HS
�b9�'A*���+�
Z*�S� ��>�+�'�:�u�
~j���rg��	ޤ�'�"�b��$KU,t@��M3���'��8�H��dK��Q1�^~
@��'�hh��Ȃ���yc�ȶ�nL��'�(���8�ԅkU��x���K�'�P8��
LAk���.��h��`!�'��j��^+q����dgN^�4�8�'`�A���{��e񠝉P��h�'=b����b��%
Q�]�LRFD��'���Z&�@G(TK���G� �
�'�|�����<�8� #�P�r���'���5� [�p�oQ
	?Ҩ��'��iD�������E��t��'���hAe�0{A�]�@!��s�"O� ��it�̮w�X#��U�i���p'"O<���F]�h�H����E�)�
#�"O�H2�� &�~ŃW%I�i��8��"Oּ�Q~AZ��A]��M{�"O2`����;�e���<?v&��"Oq@
,0�H���9���r#"Op���h�R��%͜A�X�4"O�bdm��.�n :��¥w|N	sa"Oȅ����~8ȡA1��q�A��"O��S�R�@Ъ�����! X��I�"O�u� �0f�Z=�ꗆe�
pb"O���G&ɶc;���J��t��<��"O�Q�ggd\��(ң=�zm�"OL1���>V���Є�D�bΦpa"O�lS�m��?����W�`�
��"OPy��7	r,P���"�xʆ"O`�������X�=��Y��"OT�ڥ"�*\xi�� g{�,+c"OP�Pq�C�F.6�Z'��^���i'"O�����<O��Ex&�Z�Cy(U˅"O������z��鳒�!<O`�Q"ON���O'Fp����Ȥ[6�-XP"OJ0ˁb�>(��ظE)��T��U��"O�Ȁ�+��*�*%ZI��w���R"O�	
���R��D������c�"O���!ڸ��q*�ǋ�`����"O�䂐�@z�܌���K#����"O0��"��(Ј�j0-º� T"Obh�r�.+�0C����,E�̹q"O�S���|ء�&�$=�}X "O��R�?��[a`��/:� �"O<�;� �=��4�q�_�&��"O�XǤT�t�\A9E�ǒy�혰"O���N� /�0IA%G�u�Yv"O*c�&�t���r�B�T	� �"Oe��!�$9t��f�_�"�|���"OR`rv#LHH�I�i�4B�pLQu"Oڽ���� ^��E	�~�p��"O��AG
�>�>d��g��� �"OB����[�P��d� fU �=�"ONI,,��"Q�**a�*[�!�d�7:�d�V�Q�~�6����T�D�!�Z�A�ܵ��m�	E�bO��!�d��l2��#+�2 :�`��� �!���46(���J&P�y����	W�!��P�o�vMZ�B�|��1���!�C>^�X���{��=��얖o�!�ă�<ۼ�2f���I0=�JD�e!���(A�^� 2�Z�F�l�K��A��!��;wA�\�ש,H�� b�@5!�ϓ(����m�09�P`˽q!�D@�Gl���]�O��`g�1m�!���r5a%+°L{��1�Ơz�!�D
�;@X���N,�[���Q!�$O��$����b�ڠGX�,a!�f� ��X�~_�mA&@�$!�D���l5�#�JW���q���>!��/zV��I��mSԂլ��u!��^�rh����=q��sDMZ�Z�!��5Rz"@�����6DJ�Z
&�!�Ԅ8j  �d'�4D���F�!�$];��!4M�p���Sc�V$G�!����5A&O�R)>=q0$�!�d�6tF�cB�;r�Yc��j!�� �$c D�u�ʌ@�R�5/f�s"ObP�����C"��:P���*�0�`�"O�9�J��:�H�;��&U�
5�P"O���^XI�����9��"O��X&�֕F]�Dm��`=�"O�ŲEK�6=a~ɲ���!J�{�"O4\ɒ��-+V!��%g�#"O�%c�Òr di�Hج<|��"O�� �鄌uܘ�'��O�|�"O�t�/�R<p8���9�@��"O��QV�D�*>�h���"����"O�|Cq
�1�t��$i	(P�zM�2"O��Ы��)�q�Gǉ�SbF��"OB���  �   \   Ĵ���	��Z�v�G�4P��(3��H��R�
O�ظ2a$?�K&����4`��b�wa��2�� l�B��"#^
�7��Ԧ={�4C�2���:�'��&��(� ��8 �� �L6xT��B��v�`Od��� 0�O��_=	`�@�NC�^�p��Fꋈ	�,ё�\Cy®A�����tgI�����)\j�)�6�����W�8=F�k�΀*d�`g�,}�z1s���<��$។A�T)O`��D�ֆ ��T�ˬS���3Ҫ]!x3��� �x2��w�b�����$��'j���'�n�"�<bΪ!��EBdiBL��P��r�O-P�Q�(��|b�ҦL�x�@�Ѳ.�`�����yOOX�'f�FxB�7� \�%BQV4�p��7��#<��-�a�"� �,i���6H"rlH]��d�O�mh��?�'+���f^.D���������Rݴk^,#<	u-4�j�P���mU�}�ƜJW��Yg��q�Q�F��#<��h!?� �`�J՚��>\�����`�Gy�dVD�'Z�0�?�R-��	�sݏ���Ќ�Qլ#<�0J%-��d}50!X��[��3�ߌ�1O�#��D�!��Y��т&����h�@�>
��@��6Ŋ#<y�F'�I��
^9���;� JDb�S��'���ӯO"�y"�(_�1�|aa���y�×�#z��0c��;*���Dj����/P��r�|⍗> �@J<Q�*.rcJ%
�G �?H��MW�3���rTf�e�	h1r�C��4�Ie꼼��U9%��Řu�Ȝ�c��XB��;��  �$��U�<��C>A�qt�V5��|hG�g�<�@cE�0a��+z�8w+�K�<qTaU�D��p�lФ_z�����G�<a�'־P�b-�T�P>�(�@�G�<a 
(@͒�z .��?
��1�j�n�<��&=lH i�bI9B�!���n�<Ir�ƛ4�̈@���!p�!@i�<���Ÿi]L�#J�P}�����b�<IRB��"�!��	�Ĩ�wD�^�<���8p 4�J�u�N�Cv��Z�<� E�d�Ҏ��!`�� y��RT"O�p[ŧ�޼A�4�@m�^\��"OX��H �2!z�� � z@dxҔ"OF$�U�ܳ3�D���h�7|�jp"O�;� \\�01�G�	���9"O�	)����,-�p����R��A"O���f$�>Bx�)���	��"O�   �  o  �  �  f%  .  K4  �:  �@  G  WM  �S  �Y  `  _f  �l  �r  (y  i  ��  ��  3�  v�  ��  ��  x�  �  �  �  ��  +�  ��  ��  4�  (�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;����i`9"�ˁl�$@��- G��D��O��2�	!0L�Qd�*��PZg"OJ�R������qE����Li�"O@ӥg$x�|���ֱE{�Q�"O��"W����i��ۇI<���"O4)遪@7��P�����z:�!Y"O6�#�`��U�|����%(@"O��J�΅-����		���	շi�hC�I�(���Q7n׭A)�� ���G22B�	�{n@ 8%�@��j�;(��!@�C�	�/���#�"[���@(K�c�E{��� &a����k)�
Da��>�~���"O����<A)
H�B�%`��i�w"O̕(K*$r�"�d̩�XС�"O� �fn�-V�&�
C$M&0��RT"O���T�'7_�����߇ke:%��"O\6�&un���'��V��
��6D��xr�@�I�H�j�O
<��x��"4�	}���Oi�s��Ki����Q�7
XJ�'��|A���{JT���5�
�b�'^d	�u�Y<��k��}e>e[
�'*j�� ��,3`��{�[u�m�ش�Px�E7Q�I�T�[�\���)ȫ��=���|�!�-%Z�xf�@�N��P�d���y�E�0P�ܐ��K(L���;R����'cў�Oz4�c�Z>��H
�B�Pu����'���e	ݬG�.� ��>P���'� ؐe
T	v� p��_�R;�'��<��ǔ&�v*�)T�AL���#��;"� JC@�X��L9,0�@��"O�u��"FKT�D� �ԧ}�h$""O�h"'�;Hs�Sdd��op���'Vў"~��&L(
m��nS;#g���¡X��y�W�z�B)�֡ڞ$�.�������yH�jT��ߑ1�%R���0�yFR�5X��]�$��,���y�)�6{���Fj\9N9bT���X6�yb��@f�\�Z�RC�߀�y"��KN<�P�O��+J� ����0<Q����)+TX�i�)�d7�����Q�]�!�E�8���P�	�<F٢6쓃$֢=E��'-����@,S�b��7��`H$z�'���/�r� #TfΞfE8yK��?	� ��3��.BD3v�/�>����H�MY�قG�1c?zib�e�8ʒB�$q�zA�''�m�L�?J�|��O�"~J���/�  �@�ӫ�"J�I^I�<	e�)�8D�A���MM\�	PdC�'��yr,G������C&�Zr�E��y2]%B�F��S.˚<�`�Z⡐�y�����������"1��أQ� >�O	�'NQ>9�0װk��18�)+u~mɧ!$D�����p#ȰR(�<=ެ��Se�hO�Sb�)�Ma�
R	��Ԡ�LK2�U��nNZxB��nՖ` ��5�hd��O*]
R�Ӵ �ia�F�GbJq���D���,i�i��9+��PC����!�M1Yl�)rfA�L�L=�H]�!��	4��a��,ۊ_C�ecwf�<{o!��B��j�S�ȧf#�p�$F݌5X�^�h�<E��4O���"$%U8���Ýzsb��ȓ]�~�bh��J��1�SZ��}�ȓ
V���`ǔ1J	9e�O.�8e��I�
�v�R��Tي@M҄�����ޔ�y��=R1��Q�>�<$��8�y�n�e�Js�"G��h 1aU"�y�d���Y��)9&�]��2�y��� ��U$�.;�虹#A��yˇK7`˱��_�p����yRF�&s�L�X���N��y�6eǍ�yD��{˒��F��� z|:����y"A�;p!��`�VΌ���'�۰<���̵~����A3?��!
�����!�Dә~�X���L�.�xIyVQ�c�!��\���8ׁ �<�.D�C˅�z!�� �B���ndt� "G�T�tR�"O�LB &t��]ZP P/O#N[�"OA�Gx�����l��I,�a��"Ol�����-! �@��I&3t���"Oz��e�(o�2E��gH��1�"O5�1�+>ꂬ��L��_�e��"O`��5��#J�)�3��(�֩�"O�=�s!�c^t� S)�q�Dɂ"O����v�n�Kc�������"O1:3���,8�u�@�S1�ّ�"O�xjW���4�<��1ę
*����'���8���\y��`,A�i� h��3D���i1)��K׋Jd��TR"G/�nӺ#<�}�PB�d��Ђ҅�F��a]@�<��k`����q�]x�t����Q�'��yrj9
�ہ�ĕI��ڥ%�(�yں�v]+P�J vM�8����y¨�Q���
�>k_ ����ybD٬Z���@gG1cpuZ�ɔ�y�m����J��@6k�`:'˟)�y򣀿��U�F�ZmyrP�L��yBf��=~���cV-c�4-�F�&�y"�m�11p �)^[.�ň϶�y��K/�9Jpd�JЬ��)��yB./M��}���2F���# ��y-�*�	��7�������y���8E�Er3���'����D��yB��k�<��w�"��ӬC4�y"��/7X�RD�j�J-�r��y�7U��)&̒?s��2L^-�yR�H��U���X�W�$�h#S��yR"�D6�E�&~��E���y�L��14��2咿"7D���
�7�y"GE�� �#��.J�Q�K��yrN�9Y��:ebR���U8!��yRE�]�}Y�!~J� :����yr��=	NI�u�D�!�8ʗ��4�yHI6�zb!�	���Y ��7�yR��r�V�����
>��H���y2��" ��ܒ��ԛ"p�����yR�
!J�f�Y��	�\IҊ�0�y���f��2L�
㔍k��A��y�F�:sx��+�����siC �yҊؑ��M�2�� r�X �m�yb�5a�e���X�.��*��y���q�| :�腼9ْ� ��yBEϺI��Ȉ&�֗8<�@�F<�y���(H#�X�z?(�zP�Z�y��(E�0%V�K�C.�21ې�yb�D�Q&�۷��8J&u���)�y�x�X��膛9����
�ybE�f���%�h΀����y�k?i�̺Qώ>=������yR/
g��@z�c�!e�(�]1� B��.O������tm��җ+"RB�I�~5�wHP�Y ��V�V�NUB�ɁRRͻ׆�"*�T&¿U�C�ɳ(��LPU�S��Y�_J��C�	�tx�QB̗A��c3bX/)��C�I*aC�]��Fߒs��5Hv}FB䉀5�����i~k�ꔟqQjB��K%{�`�>m墵�B`_(/ݤB���A`�.O��F�
���3�xB�I%�!+��X�Fi<���Έ,,$(C�)� J�c�O;}n-�$�N8E��i!"O��z@��t�N'@K�h��q ""O�*3쓳1�	�C)�2�@�9�"O6tA�͕�)�A�'>�=��"O �0"�Mb�%��8[y���'%�'���'$��'e��'s��')ґ��  Tz��# ��vX�4'�'��'���'w��'e��'^��'*���)߁9]N�����<V�QW�'���'���'o��'c��'"�'�|�Y�Η0{���6
��j � ��'���e�i%��'�R�'���'f��?t�X�(s,N9j2S�@���'���'��'b�'���'�b�'݀<
�^�Aڰ����Ɓt�"�b��'cr�'CB�'�b�'���'�2�'m�4��lX��̴,��(�K�7�"�'��'���'���'�R�'���-��� �ϕ)��t������'?��'���'�B�'���'�RMY����)�.P��<i��>=�b�'`��'>��'���'F�'��J E+*0�d#Ӯm������E�B�'+b�'�R�'1�'{"�'����4NyÄ�@5�d���X�)�'��'O��'tb�'�'#�g�43l��&�"b�2���VP��'v��'xr�')��' r�'Z"��&xܥ�̃�kV|u�M�Xr�'��'��'��'�T6��O���XT����,X�b�jq�#�öy��q�'@�Y�b>���&�G,��t�N��K����a�*A2z���Oz-oD��|��?Ac@T/T,�«7?G��s���?���~^��ܴ��$v>�������/O������R7F��`��� D b����fy�퓜er8�ʖ(H5΀Q�m��/g��ܴF�&M�<�����h��Κ� �\ܳW��+2g�Y{���r�,���O �	u}���$��b��f1O0�;wF�/����$�%Z�����<Ox扽�?�U-/��|��)���8���A3�E��F�sC����d*��֦͚�l"�!n'&��7��~���"�%f��?Y5R����۟�͓��D�6K�PXQG��A����;���xI��v�c>yA��'�����e}rӒ�	��n\�r#�)G�l-�'����"~�*�f��$���p��iu���Bg����4��x�'h�7�-�i>�!����������5j�q�����|�I�h��en�Z~25���ӀRg�9�-��e�'� UP�y�'�8�a�eB�(� �K��\I�n�r�'�9�gF�o]�\Z��D�h����L@�Upz(y�d�<bti�_9k�,t9�%��}x���A�|��E�GOG�I
��B�#�/JJv� ���}�Y�b��1~JZ(�g�(Uy8���&brM�f&�9f��a����i�H���?bYf��U�ĉ�R�#$�8R�N Ǣ�b��p��ʧ�0>�FF.rx!!�ω�N��}Za��v�<i���".��b�K�*z&��tl�p�R�c��,��`���A�Б���#3
�aZ�N� Rv<��o� iz��ӻLM��s�E�Rx$)��mj�#1����$��N�6�:b�ح`"Გ	�Q��A�톢5����	��Z�R���麰k���{	lXS㫅p���Cg��-l8ېn��|L�����2D���q�� 䜝��������C�	"wTLڇG��\i�}�烏7Z�B�	2U�-#T�
�(�1#�'&T�B䉷Q>�0���óU|��{�(��pE�B�	�G�����1l� �Kܔ!#�C�I�x�h�E.���A`$hբ�`C��2}��)�+P-O�P��1O,n�dC䉻SXj����'�qb�ΫN��B䉣'-:��b
���l�-֦B�ɲN;��$(C،�FN8}�B� NI����"��iO��DB�	>O�ꉙ&�_�=d�H�B�nv.B䉼�L5� Oއ&�ݘS�U7m�C���hE�s��4��4[pH	�C�	"` t�JG%[=
��(�&�-<C䉎6�b����H��s6͕5H� C�I!]�2����Q.�Sb�֓2RB�	��l��ȗ/4�	�֚��C�B5d}�(�7]3h	;���&D�C��	a�\ڱm½[r ֈ�Y)�B�	�Yˊ��A�u	˷�F�A`�B�ɚ[��U�N��c=Q��ȅ�C�	,��l؅�ɣR�4� @E���B�ɾ^Qf��S��&|�85�!� f�B�)� �0c4�Д�f���iL'	��y��"O�B��G� &��Jo�����"O��SV��nN�"��o=z5��"O�e+��՛ ���"C�ҝ 7R=�
�'�j9Эځ�0�w��YBpi�'���c�����$$5	0�Q�'��c��p��2IF�6����'N�t� �
#g��9���	2���
��m��u�4�ТU;�a��G�{�h�rg�S��d���!��e�|�*b'��|7�>�VrqZ|RB���b��(�O�rXaӮ�;m�F�i��%c �	�'p���1?MX�$E�Uz�u�'-����P�e�ReZ�OI7 �"r�C���,��Mָ~�|Њ���n�<Q�eD�s�B@a�DĖq�*�h��M	u�F;�'f�Dm�R��ܕ��O��H�0t�b��W��_��� @�'�J"A� =��iC��W�jX'LԀ9���h�+[�v�*sѡ���0>��FE�5��\�E�ߡk�tp���I_�'��Slz`�s�� ]�r�{�?���8��W�i:�s4؁yq"O��8uGY�V�c`E�}��ƾi'�)�˚� ��铤�Б=Q��q�t��5�!�$����4LV 6������ͩ�y�&2��M�d��Y�25��O�!��`#��lӘmq2F�F��h7\?M��:p0Ġ�����5�Ã�a~��Q+�Ԁ�Ղ�.5t�����+�����AZ�Y���PG�{����IE��EC�+U7��87�D�*#>	��Ù(�|�(�NͱYgF�r�P?q��/X�؝���4JzXh�&&D����"w%�(�&D���ti$Ji�,pS��/�4�B��Y�"��	���O�e6���(����3g$G$;N!�d��� �( *�sNx��ϲ>�&�����e:g��B/0�[ҏ,Fx�f�5"iT��e� \ۄH��B?�0?�T���ws��0��.���D��,}����ɬLs<��%H
�Ta}"��5>z���ɔTt�2C.�)ֈOD����W/1B<����=��d�Oܖ�H�a��~1Ն߇����'�rD+	&K
j9�s�^
u1�xڜ'4�a�����~G�RK��7�?1�#�Q	@��l��O�<���)0D�$�V���rP�@�bX��3"$�<�e̫!�2�	3Ƙ��0<�&���v�lK ��\��q� �pX���	% YD�Ҧ�ũ#N��84*�	Y��
���-_^��#��#��\~��u�6���)$�LDz�nR�Q��X��)�P��kpX4 8z�b�A�/!!�D�6��h���4#Z�#Ʈݯ	���M>v�9�=E�ܴWz��	�0sp�x����4��I�ȓ	�TI#g��\o`9�������'���x�'6��Q���Fς*6�B�q�춄��6OT��u�W�8��dQc�.=���"Or����/D�4!�΃&N)#��	�-���ق��*�:]����-m�r�k���=�B�I�jm.h��˺? ���M��6��%M3�a[���s�
cd�"�:EŻgD:���"O���@8HQ�)�LI�Y��_���D�
��e��ɝG��|ᒆ\�d]| �� #�$���� c $�{�|�ܕ�#��� �$��Q����B�	�V��a�� ^�D��pQg�R�V��'	���N�L`�AF���6�(� 1\q�� �j�Ӣ"O�ib��]F}�pTb�2��]�0�'o��R��J �??�Ϙ'��i���u�,�1�Ewd�0H�'4�k�GW�v��hP :nZ.|�rDT	%�t�4\�]���''�I���3s�jq�#� 3b��	�-E���R����uj�$I�V�b-L�!�4���ڒ\C�L+�'��0Up\ɲa�ffVQ"�O๐a�Ty�f �lo��D��c�0q� ܀��� ��i
���+�ymE:g{@��K�C0�u�vBC�����=�r����S���~�<Q��-0��;���"��L��) ^<Q�ˍF �0���#1��Qc���V²�oZyy��
�\��N���DQ=	ANa��\m �ej0.�axrS�/v�nԑ� Hp�L���d#'��U��B �i����	#�O�p�GQ�z̪G_{J$d����Q'����3|
�E¬O�+�L�?m�tM�^�u��fȨA��V�*D��$��M+PE��8���!Jh��۰
E�j����d��?�Q������Q:`�ᝡ[W��yf��[U�R����J���&7��ř�hq閼i���I{���:7�
n]�4��'q�n#<i!�2OW��S`'N�}��$�s�'&�x��e�"�M���r81i%�'/vQ�s�ʵx0 ��j�D�\t��j�}�]9�p������9Hq�AOAa�>�D��/R@�!nZ1TV����������<ͧpE����0����� �(\!��$�\�3�CD�@)9@�3'��@F�3�D��X�p�s8O��e���{���y7I-R���Q%BC[�����!���?a6g�$�58 �X�ZH�!�ɢ^v��fM�C���Y��c�V��S�H��#<�3���MH��� ;{��!R��D�'Ul@�$w��y���/�I@�~S��*viعzT��y�CKc&TE�3m�̦9S�Zt� I�cز\Y�����X8<&����ȧ>��L�-,D�dD����~��|��iA6;�J��r������P��K�<��b%S
� c�^������Q@5=O�t��IH~����y��W�p��:���,Nf�Y"�G����?���ˏ~a4�`�b:�����gSI��lB@G�)�~��'��84� "<�Q&��S*H��Y$�X�C�$�Z�'�t�PE*�56H"0
�"������h;l-�d�P�v�b2m�.]�	�m.��Dǃ��y��'S�s��а`�*m��I��B��%�Th��1��O��PĀ(�?�:`c��
�@�!�޴F7���#;0;��Ն
���Lip��<�����t���g��CEm՞b~\�jc�ߥD�B�h!�EB؟�J��ʊ}H
�[�σe�Q��8{I�����5��=Z�!�O��
Sj� 
���/����I��M��и<��"T��~ң�B;7��	�/ �Zy@	��M�<y #˾W����ə���;���q�;v��9p��쨟�hE�_�s�Y��S j����"OT8�
Q�q�<��Q�_K�m��C��������h��$��j��mK�ΆX�$a�� ��;�!�$�8R�;Y#�80f�¶)�"m ��`��1�'�VXڰX�5aJ\{$ W��Zۓ+�"�"1+�$� <�R��5�jl���VJ:!�$���x|�"�fX��*��ұO�H�-��|
��E��'��R��!�oػuV�t��j�ykP-y�0�F!�I��jX�41�������h��$^�Ԛ��f�Q�P���j��E�!�D  y�腡(U�� z`j�:4��	� )ҡ�
�>?B�	g`N;hGr� ��pӦ9�1M#t6O���F�
[3��c���FP�I�T"O6L+�KX�w��ع��6�H�J��I.��ɉ�鍮1��1{�cϐCP|� �*ӈK]!�B/AyˇNɼ� ����g��(X9Pb�"~n�2?�R��RF��py�	���72��C�ɻc*�K�h�R�L�"t,�^���{0�1a.-|O�Ԣqb�;:ԑ׆?Sۈx�7�'&��c���M��O�>HL
@i\�����vn�<�ä�4�&��"oI�qLnpJ���C�'o�bTD��H��� �H;��R�*�	eb��;U"O�H�fb�)v��\b	'J��p�i^��2�"�u�S��M�b��@^�,����T�L�h��x�<��`^��p��b�Z�Y��l�s}��W%k���ė�OI8<S��+@@�3wo�>h�a}b��v扞)b��
M�S�\<2��U�B�	�.�Bp�Z=_�p˧ �%+�#=YeU'�?��v�]5[u��`%�<��b�8D���:7����0���.9���w�@[��M�S��M{����&f�LȐ�Ӛ�4����n�<3�����%p�F�%CȂ�xƯ�k}�'��V����M�P6|}����}U���c,�dK�}b$�=�~��Y�d��G�Ҧ}��@2�y
� vq��rM*L�����Z��`�"O1���2T��(r�Z4f��Y��"O$p���E�6t�P�B-�l�#q"O��aW����]Ѥ�]2ZtF�aV"O.�`æ�(x�:h�,�fX9Ѥ"OPI�7
�!e�|���NHp���"O䝛ǭ�mT�;h�4[�8e��"O�,��јs��|Y�ś>ʸH`"O�Y�q��,[,�HG���tv"O�a����dal���D������"O��SH�;�~i@�f����'���R�XVh���gP�D��L��'Px��a�c0���g�/l�ER�'�>�J����tٙ�!�$���
�'G�=5/�9�eK�7
0k�']�=kd&3`�QEA�&e���'��:'D[-v���H.
t���'b`X�r�,<FX�ABړU8Z!��'����Q�N��I��h��_!pt�
�'XЈ�&�/%Ҋ�QHɯW( ���'�����e��I`c�JH�u��'��4���� u�Θ�d+K:	��'30�7'�).���^�1Q�}h�'�<��5�ӞB�"�x��-xR6"Oᓑș�r�kFڡ�i�"O��܍nix̉1�|`#a"O6-S&*ə0x`����?`�PI%"O qx���
e�	1��;W�EZ "Oڅ�׬�7W�����6U�%c�"O� R�7�@�B�n��،"O���n�6�4��-ۉ>�b�	r"O���I_�4��]�m� =�ڰٗ"O 
$!��*hj��H�S3V��"O�=�X���Z$Y���3"O�A��E�/��:((n�Zq"OT�@w���w�-p�X��bM>0X!��@6�P���-��՘c��+bI!��^�C�F���
�]��в	�!�d�3bК�S`bX43�$|��͊!�Ď= p��T���g��P����!��I����+pj�w�`EaLZ0g(!�GP����"R<fiT�K�(��&!����6��$Ό/��4a�>)�!�B/(O��k`�������!�_��P�h��Pd�t ��Ь/!�d��	e�M��-^�>S�8zvj�	�!��O3Ծ�����8FԀ��K�-	!�!��\��	֎>���H>M�!�Z({T��:��ˤ(� 2�A�!�dQ�o.���ݞ<=T���d���!��/i-�uP�˖)�Z(J��W�!��Bs^v��%/	+#��r��k�!���$툴�De�2#&��5j��r�!��& �}�3딓F����&�,�!��ڞRb�쑖�H(t�`����`!��+_�@��[�Fgd��CU�6�!���0�2`��a�8y閉1c !�$X�*��H�s�_�Pr�U�� �r!�d^]LPR%��x�b#�.��?�!�ė%)N:���%H:�|�U@� 5!򄃮o:Μ�@`�2G��~�\�'����O=&��&�I����'}�	��aU8C�@�xF�{��%��"O&U�����G�l*P,�#* �A"O� DMh�F�Z`i(���J�I�@"O�p%ʌl��M��F[��1"O$��-�*$�Z�h�)c?hux"Oh0*�@_�<�f��塎�6Re�#"O\��b�-{���Ч��G��Ћ5"O,�S��T<4\�y! ǻK�D��&"Oڅ� �T|@�/�#Y��l�u"O�KcV�ml�`�:/��4Z�"O��q�� �ƕ0��vyޔ�"O@#S�Ϩ�@)��>c=���"O�p(F��u>�IA���;|4�"O�xе"��+�0��ُ�Э��"O�}�5��J�NHxg▣a즜��"O"4�E�*Q�F��� ���	�"O�Aw�V�f�6�P�+�����"O��@&��9���@��b�(bF"O� ���Y�n�  ۨ=VJQ�!"O�y1�gT�cT�� �v>,��"O@9zƣ�aTP�����Œ7"O��V�S�x�z�BE��4��p�"OJ����b�N�'+�0�┚�"Oʄ�����b�t�gi
�z�nQS&"O��M���R��W���|�,P�"O�m�gn?|���B䇷l��p"O ����7��fC�0i�x(��"O�$2��֤kNܱ�� Kh�qkA"OZ��.�9혭�� N�]:c�"O29Q'�]�Xy�E�`5�"Oxd������$D����<}p\8"OؚU�-�{W䒎6|v���"O|@rw��!6��3CS�o����g"O�)���0\�ɨ�O�]ap"O,�z��ܦU��,��ȋ{�n���"OB�x��E3 Q��U����`"O��R�G.i������+0�5��"O�����/%#�x@���),<~���"O���t'�>!\ ��9a�ۗ"Or��V�E�����6/��"O�A���T"h�q#�6�%��"O�����E1#!^�7�fp"�"O��;���iQ�M`a�ղP@q"Oza�`�W��D˂�F�S�8�6"O�5#�6��4Hb'�=?D��"O����J�Z��Ʒp>�l@"OȅB4�ҍL"�I� ֝8�T�"Ol�%F�L�����nS� p� u"O��ҠL2v�<xJ0K��$<̳@"O�!��K-J/��b�)N P�r"O����d@���IxǇ�>' #"O�H"4iԚ.�0�2�fC�r��`�Q"OJ	c�ˏ����p�[-lԎ�h�"O*�S1�ŧL�~ �bؗ3��=C�"Ox1��O��_{.P���ڴt��ѻ"O,8�`�XP�C'�
�g���"OR͋�B�>x��!��4�f���'-���ԮS+ �p��4ɆQo�I�' �5p�G&+�4�d- }�tB�'� �jc�݁W,}�����x�lu3�'�@�&�#a�Լ9$f�wF2qZ�'�t���ہ ��Pc�ov�`���'���C̋*�2Xin�oPT\��'�xy�C,]6.�R)�qf�3?����'z�x:RL�7'�i�g(Ķ&'����'C.�r�B�tyw`�i��a��� BE��N��m^74˖��*O�5ӥ�ˇ[K���`خd\<̩�'�zႄ��<�h'�T'[e�mb�'��-zC�E�k�d8�VĘ�_Rk
�'o��R�^1G�6\�&��R��'M�@+uE��D���&�"p!
�' �)�M�7Z�d�X�h FŶ��'������=m�R5	�/r&���	�'�8��Ӯg�p�P�_�kJ2��
�' �=��A��va���éQ��dP�'�B��ٝM*�$2`B��(��'_"��d�ֿ#p�t�'�^��Yi�'pXqї��$N�`����V�@�'<���,�"\�rؓ ڐ-!�=��'4\<��g
�DɈ��)��OoD�P�'�$����\�K��M��:����'\\����O��=��$T��n��'ݒ�y����R���5@���!�'#N�j�n�O��@��,�rd��'�t�c�S�QD�A��L�V��P�'���@EO��Q��U`�K�x��
�'A��
B���B垭V] ��'ӆPZ2�}E�I�L��\="	�'�x���׬�by�en6����'���"���(I���'�Hi�	�'K�-�e��ra��
 @j��0	�'O����N�T��C��7@ eA�'.���tG�3.?y�딛�uS�'�*�A�A#y�)'��:~�"}��' �T��ܶ	`���^�*1.m�	�'S<�Q��'@n(���l@�5B�'�����L�#ˎͺ@L c՘<`�'���S�ʪ�,�{`	Y^in�8�'Nb���䛔L�@���n�2[�2�'I���+}C>�z0f�)kR�d��'�­,�=��i�" PX�<�'�� 	�M-}��	��^.5ʶu��'{��AS��,�LY Ύ7��t�'H�i«��z�V 1�x���'���˕ޗ6(��s�V&?fF�9�'���#Gʘ:�L�Ci2�\�H�'�Ґ�dh4zp��R�"U��I��'��Re��M�p!u��< :
�'�5S�E=V���C�	 �l]Y	�'��5�D�5_,p��ʓ�4)	�'i���� �G�8�X"+�:]Ĉ��'� TY��+f�v\�Q�^�N�D��'�YzVY_I��*���
}��u��'��C4-A�B�h�� �y�����'���۱M��.���RIP6�a1�'�d�Z#��?SH� ��U3�4dY�'ӊ���W`�<��1�N_����'%���@�P�H��8�ʍjR���'�hyxSo�}8���ޔo�8��'I�9C��V�M�4q#Ю2���'�l������GhJ��l�&�1��'5,���@�0�`�afFޕ[�� �'&�$�S��T�☀��S:)O`h!�'y�##�t���@F���W� �'1��b�-��%0A1㤆5W�̹��'�����o.%������6K�<��'���A������K�a�>C�����'|�Q��վI8�ae-Q�
�'��P*��L�B�ȯ&Xf���ô�y
� ��
�J�6O<<�A�30�qD"O�EK@KЊtn��Y6-H�X��\� "On���R�XDt*2L��(R�	0�"O�]�b�G�rEN	׫�>8���"O�x�B@�1o��P#�ѫr�"03�"On�'�#rpڅ�f�˿k���c4"O���F���:4��ɐ2�dq/�!���(x֌,p2
	obuxq�2X�!�ē.U��H�B��m(�ቄoS�B!��P9K�@��V�Q^z�Y$!�� �!��%g�uJ��K�`��,a2��!�DP3J� �*N
{�X�BnP1?�!�$�\�i��]�}�8�ycك`�!���Z9��)�<(�V�#F�[�!��ijzY�!�� �̈藠͌p!�$Ɲa� (���цu�`����מA'!�C4�y�2�߲!��A�r��-w!��S!}��$6 H��B,Rƍ�_!�ڬx��A�r@P�%w��y���F�!��A2`Y�C\WR<(ᩉ�_�!�L��yv�ěHr��v�!�����&�ϞkB4��2)>Q�!�d�"�����yR���.����'��jM� ��]9aC���@�c�'8�H��'Ҽn�"�sS��*}8xz�'�D�rSȝw��I��@�HiJ���'�Cgbճ&V�AJ�d�j��i!�'��i���7~��Ќ�?d��б�'#����>�	�$�ܴZ7YR�'�jL����Hj��g����'J�b"+K�S��!;�*ѿb�^��'*vaB�?Q�tbwѨ�F��
�'jᘰ�ƥhwh���-ƢW�t��'ƪ	��ՇOph�+g��$TL�1��';��Qo@�+�)����"�p��']�x�"kQ�t�2Mz����-�3�'�*\+���'��ؚ�d	r�40�'{28��"[,�[f)F ~�A
�'�4�aᇅ+�����h����'�l�q��V�P��SbM�(!��'�:@3Ƈ�C+ ��H��X�1��'�Y`�.\rh���.U�����'��T��LA
K:�r�M�d���'�"}� m��BP] $�I;pmY�'�$��nx����K�O���
�'��Y�gB�C�l8�c�:��
�'��C���rM����0�	�'W�ܨ0M'"|mH��� K���'\>e�W�O>:�X0� !q��[�'hЙsU ��@�*]�".U h�d���'�sw�va�염}c�a{�NP9�y��UL<�3�O
o�52G���y����?BhP�׬�gc���3�y�"=�(��Ja$��!DD1�yb;�Ht��0%p�\�A��6�y�ϋX���+u��R�L5Z�H��y҄�N���$��*K�-���Y�y"��<�NL��!:�)�v/W��yr�	Ln��̈́(:1Z&+�yb��$x� �@�6�����ͭ�y� �?|%(ŌI��M�#LL��y�Ç'V9��� >5��e���8�yb�I�nW�3�倒1�5�����yROO1;}��8BΝ�#��ٴjϛ�y
� ��1c�*E�L����(I'��$"ON�Qp'�` ���m�}08IJ�"O�*�H��/� 詆Ʉ.�%	�"Ol�8�A�<M�6��̊�>Jr�rA"OxA�N�"5>`U��k�e�lp�"O
P���:>�6eY�I@'U�8kd"O����y������` �u�"O�h�Ϣf��p�Dr�2-��"O�]ɡ���p3d��k�b �e"O�I�Q��1��Iwb0v���"O�y�J�!R� �A!CW�zeX��"O�p
��Їc�c���tN�(�4"O�58�E����ī
m/eK�"Oچ�ĕ!��E��#B&"��h"O>e��Q�Z�zQ�7���"O�)@'�w�81C���+���"O2�hgFX#���w��"�P���"O�9�T��`�N ���:;�
4iP"Obe�		dAr�@#'�U+p�#"ONX�(͚-�`	�L*-~�l!3"Ov�z§�R�vx�+L�v\*Xt"O�Q���r4�K�L �p���T"O���S������K��W��]�`"O��p�B�,<�b�ː���`��"O���C�O�$�k�ʖ�0%�ݪT"O����ڠxL�@�ƒ$H�=;!"O���l��%�Τ�Q�}��1��"On��玆*�d�Y%i��V�����"O�P�U
�VL(qHZ?>����a"O6a��B�c��܈�f��j,��"O� K��Y���j��8��Q""OF`��!�5:�� �]�'�B� "Om	��D4 8J�e � BiH��g"OzȔ��
�hC�O�d�`"O�U{��WJ�&=��-KZP��˷"OEhE٤?����g�ڃ"�� 3"O�u�r�N� %�eA$q�]��"O8g�ڨ
b�q���zb�9{!"O2�km0��Y��Z�ư��"OTkBl�"5et9+S퐃=�h��"O�ٻs� ���i�̏8����"O6�2��ڸ%}��+^��T�Y�<A�.J����&�$m�Ұ���PS�<����K�z2�Fzn��&�X�<A0�V
����N�����W�Y_�<�cu�8`�힀$��-�	�t�<0NT�sW��`�#ٗ7�(�t�Fp�<qv�^4I������^T�񣤉V�<ф�jCr�X3G�<'�xM)WS�<�u-݀,`l<s��6S��0#ʙO�<����̣r��>\*)�rD�<m� ���UA�?R&���aYK�<)����X:�L�AT��扙�OL�<�1'Ā��=�Q! 9%��m�A�@�<AS��	c$�x�/	 C�$dQc��V�<Y�A*6���@5�J�"����l�G�<�7 B23�|ȁ!��~'�]{��G�<!�Bi,�1	*��S�h�<�@I$t/H��S�·*�ԩ�nC|�<�.�54����E3q�����z�<�5g��|y�n�33zT�,Y_�<��e���$��� �?*\�7/[Z�<yQĞGJ��@���,<P4�"aC�V�<��I�+	g;�*P�x����7��T�<� 
�y�ĝ;t=r��0�X���q*T"OM÷C�J�*}�I��6r�}�u"O�M�WO�5�j@b�<Yad�"Oh���@D�BE+ШÔu:`��&"O(�Z)��C"cS�*"��&�y�<���E#���R�����)v�w�<AW�ڃ7V�j�����Yv�<�1�dq�IF&�~�Tц��G�<��@/06ݺ�d�m`�3�BY@�<�Fb�s @��D���
� �y�<����49΄�G>,�m�t�<��g�I�ƭs�(�t3����@�j�<�^� H��kgC�fe�4����d�<97���Uʨ�	1�BpBz0YQK�k�<�r��r�|i���=�0�ca��S�<�#�R����	;�Lġ�Ǎh�<��D6���ҔL[*��t�2�O�<�b"�6+xA2Q/'y<���a�<�A茾{�u:�K�3w�̀�h�<��i��|���(��D��(XC�A|�<i�e��:k�2�+ ���ţ�f�@�<A&�"l^�Q	vo��h�@�c��T�<�sϘ�a3�	�K��ui�����RI�<��eS�B�� �b�20<������<iR@�3d�p�p��B�)�|��Y~�<As!X��=���U:6��dK��TT�<ipf�5qJ�0êH3;frh�w/E�<����&���,M�iW&�hcJ�g�<����):�f}�$*�{�*æ�`�<)E��-~��3��A��.Ѫ�`^�<� �4���i$"F�D�W.\�<��Fsюt����#z΄�dD�Z�<��F%��P��� ��X�<�thN�jg�Ѐè�r��%3�!JZ�<����$%�<<�q�XI���C�z�<�Ҙd�������#Y�)�u�y�<AS�J�=�T� $�I�.y<��F�s�<��AWr� ��?�N���i�<�lX�;�0U)�gN.]��M�<	���l�.LS���u��b@-�J�<G�ӂi�K,o�5W�O5��C�	�)�J� :��\�5�Z`�C�I�Djh4��[�uT���g�RC�UKj��o_,YT @��(|V�B�Ɉ3j�9���B!	��ps��PB�ɨVC�ԉ�H%��p�M��$B�	w�>�Ӡ�Ƙ]hv��ă�7��B�ɑ1���e��#�F���	�+g|�B䉁&_��;3f�0y�.�HQ*�;®B�	�o���9��N������!D'!�DɲUD����)��<��`�!�D�dr|r�� �����*��!�B�uѦb�UxŲ����J�!�$S ���G�L�r��V	�!�䕉�¶��/Li\�q΂K�!�+fw��"��	T��%�N�!��I&!�����!�!�d��R�!��Z'd��ЇQ�jxdW��9�!�D�'�x C�c��[�ف�O�2?�!򤁽�䔃�6'S=8 ��!L!�D�\�khG?�샴��!��٭<dX�ڷi_m\JD��KK;:�!��|����oQ�k��-��I��!��	$U�J4���ùj3j�[�WG�!�� T�Qe�b�8�1��V�Pw"O���B�)�Шp`!ɓ����"O9�"n��7� �Bb�	l��U��"O����ֈ0ʙ*���2�X�0�"O�m˖���Ux�4�_=�[�"O ����*F��YpdN�h&~�r�"O�-�U@"|�)���� �xy�'"Ov� `M�v�`�%s�*	�"O�}���|3"-�@�8��x��"O2�% P�K5+��� `�� ��'�ĝ�E`�;(^�x�'쓀��L�'p����N�byĤGj��R\��0�'�0U{�F62���#�͈E�d�1�'}����U3m%h�p��7�p��ʓe="(iGÄ�nQ��{ �4-Ѕ�3j�R���1Ϊd�dʞ�( ��^���
�ǘ�z���`��#ֺQ�ȓ`;�����Uj��0�b���p���Z�B4��3�"�&U31P\؅����lܣ�Ɓ)p,�	9�H�ȓ^2PD���$/����������o��m��ԵSt�M�@�*��@�ȓ�*y�6�^Q6h0w#� Q��A�8�3,	]�6P�+�+��A��:�Fy1� �7��s�J�2 ��r�4�FFɆq9���@�} �ȓt��M�T"͞
T s�,Y��܄ȓ}SR\2�T��p=��׀D�0��ȓ)����V�,<2�I�Agҹ@��M���L,�G�,�R8���32+����"�K�����k�P&ml����'U����ITHz��)@70ͅȓrp��."iލ���ؠ��ȓap����]� ߒy%� ��5��Z
�&�@q�E����s��ȓrP��g��9,���p70*:.]�ȓ@{\	K��0[����'��2~d�Ɇ�B?�Aۦ�Ǣi��8�B�;xp�ȓ�
�:FN.��=�ы$r���ȓ[w�5"p��"�B	��m�Ux�x��pi�hR��^>��R�]���1�ȓW��rP��*���#6��54�¬�ȓ ����A٢F� �����H�^D�ȓYl�d��*�N��������ʓik����l�Q�|�&�6zQ�C��m�2!#�gR6L ��;�#��^*�B�	1{�,���VI�@��c�|�nB�ɝ
]�$(1�Z�,KL]�c��dB�	�Nw>��yr�kFAߛ}�B�6Hj&�2E�y��9S͛!rC�B��10��*�L�!�����Γu}VB�	(F����%Ü�~�ы���%	�B� �l5Cc�+@�2�#��*!�C䉃 ��tʍ�0�Jd����>b�C�I�>��M;�kR�:���*EoN*@�~C�	�#�b��F��1L%~S�'�*EuzC�I�UB�)�g��h�8c1j��A�>C�IhbE1���&O|-�����*C�I�Oz� W
�<eB�t��ԣ
T�B�I(aJT�;��OW�@�`���^sC䉼crJ0(2b���f/ΉMբB�<WR*�!�NP�� e�ԫH�q6�B䉅h��)D�޼Z6��eE�	�B�%{�MI����Tj��V�-IhB�)� �)�ԩ ���@��#=�bR�"O0tc�F�d�P��"E�0J���R"O����nU?Wwj�� �]�< �C"O̬��D.$��#"�qNH�G"O�H��aٲd�X��Q�Q�^g �Y"O�%�ĦԬb���*`�K�I5VQp#"ON03�o����,�6SI��"O�|B��;?~:�f@'f�@�"O��"X�*�
��`f\/S�a�0"O ��&����@�E\��"O�� �K?����OҰ� �v"O����c<.�p�L�y$�"ON��D�[�N��sьͨN�98�"OB̂$�Z\�5RW�׽,�0�"O�� �32���*�mKt�*��"O�#�M�5>��,A0%.zz!�$�
#�@HG�_�B�6+󂎲!�03������A��Bp��9L!�D�"6o��&!�<q@�����k !�d�3f�ܓ���#>@�I��
�t�!�$����IVjNb��x�d�E� �!��Z)!Q�ؗGp ���M'P!��t�&A���P�ǹV��R !򤉑�b�*� �� Ul�)�#%W!�$ō�~pل�ە7bʬ��j�?uG!�$��z�×�/M`(`w�2t!�Dх�lY�*G�v;(�s0l�+z!�&d��s���-s.����! ��!�$�02�����)�9	v��bq!�dU�@4E˖�ӱ,��E���_!�d\:	1RA*�.�&�*�K�
.W!�U�DC^8ǃݡQʄ��!��*XH!�B�`�(��큿b�RӤ��"N�!�ĈGse�J��m���X�B =l!�dd�4(ǳq�
�d�Rl!�$�:*g��櫐7Az2� ��	�S!�dY�ZϒŠ�ֶtj�P �
O�!�d��X7����b	X5��v�!�ç�ȑ񎒴���K6!�!��?#�D�r�iP/��z� �:3�!��#+6���b��&$�MKՄ�)t!��ɔ|�Ȕ��A`$@��*bu!��)[M<�1N �t%X���"5�!���	���igܕp�A${�!�
�EV��&�_�O�ܩB�f�(k!����*��@$�*0Y��G+.a!�E�u�\��-�z������ )h!�dO~�Fu�!V� |�2�bW�{�!򤞦]9���$�'`V �@�^�p!�dǣ����r&13��)�E �d:!�=����E�`��%	 E^G!�$�$CV*�)H���@ �k!�D�Ig�x��a�%`�e��K� �!��uCR,)`�\9S��8�)�!��2���ա]Eּ#V��9K�!�ݹ\=���P�ցX2~*SA�{�!�d� in�����5�����\�!�^9]�v�� �?0�	#d�[��!�R�<s��ɗ��:R�ȥBf�~�!�Đ�Bb�8�B�=��-A��-u�!��4xJ�����+}�*a�@��5(!�d�f �Gk�� h�g)��Wn!���A�����%F�>� �I!�d�	g��Y��Lr�ji�Ҩĵ<�!�� 2��u�UtU�����&>r���T"O�X!î?N�Ř&�iAt�d"O������aXưS�L��OP`@�"O)C�=�"}1�BK�C�� zE"OHU��W'"�k""��b|��[�"O�ĩ��_/$Yjp8g��bɨ5"OV�闆�*&ډg���?A �:"O�r��R<��e
�2;����"OL�
Ŭ�/<���S�	,9,q�E"Oa�T)f���I�RE J��7"OtQ ���ey<�2�'�4��"O��&Ćb��;2���y��"O�A�猉*,�� �kpع�"O*��'B�ۤ�P�O)ER@! 6"O! @Æ�;s�VJX(%"O�����*D�ݩd�;	���y�"O�$Ц��qJ��j&A Ԥ�i�"OfYHabзc�pHƊ���qL#D���Y::=葎Q�d/��2�3D�l�� jv���E��b�H4.2D�l�R�͖T��Iz
[q&9R4�.D�H�Q�J:U�D�����}$��K�+D� !&`T��<�p�^)Wxh4f7D��R$[% è=�tf�4 �,����3D���5+Ū`��S��Ӌ|���Ee3D�X�A�|������p��t�$D����$(0��Wi�6�����#D��$Y�>E�y`�l�;w�~Q	�j+D�����R9Na�Yxt��*wG\ib6G6D����M��+z�{�.�u�.-s�4D����B�1ؾLm�9���1���c�<�v�X K��9 �1>Cր9�c�<��̔}��ܘaD��<�|�T[�<�eD�6	�$��6��U��X��s�<�V�]W��D	�.y8���c�<!���9&�)��&AI ��5�Jv�<�2�ţ:¤3E!��Bښ�8��t�<a"E�Z!���bKT�~�tC�	0V ���5��b�"U�A�bl�C��?~h �j&�Vl�wM�#7�C�ɛvތ�i2�Q$ � dC ���C��:}�Hr��3n��<2��߮R``C��/+�R�s��1�Fes�o�"=�hB䉓6��]�3L�d���A@Aq4B�	!C��8�Sm���0C��B�	QӜ�兛�slT䳔��R��C�3D�ƨ��#V8u�4���E��C�	t.X�!�o<Q� ����C�5g~��h'ES2�Z�V��B�	�(K>`%4D&-yV�'�B�	�Z,�t;CJ�7H1��[B �/L�B䉐H�����^���a��`��B��;%�@I�O�M�B�)� ���B�Ik"jh{��${Ʊ��@�%�BB�}�l��ծ�.�n��F�QB�ɱrȐj/�,����P��rAA?D�`(uKS�dzډ��IE�`�o9D�p�V��aPR���h�v_x��8D���C�7�^�I�N'P�p$r!g0D��:׍�\���0���h�d�a�"D�����,|
TY�R�	� ]d����?D��1��6�J��%��!�F8�h3D�Ј�N� �����n*�p�,D�lK�/;�l�����!��a9�+D�� ���X�$�K��/@A@���"O���ǘ".a�L;V]�],�!ʃ"O~Ec�lS�4��1�	,��"O����0�� wB�Z� ��"O�D����I.�t�0���|}��"O��:�&�93�r�!���c��l"OT�ꖡKX������J2"O�ĸ��ɱl����Kݍ@B,��"O`ݛ��Ɲ_�`ۀ(�_CPY""O�8�L�?w>���&''  �"O��S��]=3���F����M��"OnA�����P_ )��Fħ>�lR�"O
\���N�ei�Y7��WpZ	�"O���AJfa�e(���Y[�q�A"Op��K=hTB%P`�!I��i�"OXy��G�z`�ٿT�^4��"O�V��J�!f��AM"	�n�<�d$ɰš�&�a0����Ho�<Q�E]4� ����G�u���j�<�P �>2O&( �[�qz<zg�Yc�<�c�
"}*�){w	
7'Ҩ+��`�<���W�nj�� A� h9fQ����g�<�a������@��v�C&��j�<1��	�^y2��K���2Efn�<Q�JB����!	�5� ��w�Si�<����1�J�e� O�
�;0o|�<�1���9e��0��ס��a�x�<9q�޻<8jty��֩R���'��v�<i��űy-l�zNC'd���x��I�<�I|�t �n�TX:��C�<y���t#	�`G�75��8S��G�<1��O�IМ$�'��'�����IB�<qUD�qD�q3�b�9
cvT���H�<��á0�h��U*Y80�\}�2C�G�<Yw��!u�5:�!K�4��˰(�o�<�G,�f��DRSN6-u�1#Q�<�­��t�69����1lGu�<�R,�%}�X�'���@;󏅾�y"k��r.��O�Q��H�qa���y�E�5X����ؔ:����I��y"�R� ���j֘b��y�#�yr�� LE��"V�ԽR,��cI5�y��%'7��`k�w
h��Ua9�yb�͜V��Չ[ ��I�2��y�޲l�8�`����dU!��̽�y�N�4��W(�nwl���C�(�yBJ@�R"���O��`.�c!L��y"��V�`h��A�ZA�@r�)�0�y��]�4��8��ɭR��Z�"/�yG��z�Q'��tt�8R�lC��y�n��E�`2� ����r,���y�AL�_����r�׉�8`(Q�
+�y����
u!�P�D��'�ޕ��^�>���a��C�`���'P��3���k������'��������=��&G�X��d�
�'����H�9�QX,�;��
�'
BQ�Vb�
Hh��	(&�PI
�'5L��s�/|�*�	Ӄ�$#�P�	�'9�y"q�L��~A�ʂm�Ђ	�'���2�] �ư ס��j6����'��A���)Z�� !�̘ь��'�a�Q���P�eѳn�Y�'�� pր��qL�I� I#��r��� ��v�=SnVxI��B�f_n]�T"O8�څ�2r�����cyf��"OR�f�4j6W���(h�U�O�<Y���4s�L�;���DE���YH�<$��G��H�cBйar=�C�<��S� [��A%�U[,��� g�<i���`aV ���  NN��z�<���0\Y�iP!Ȼs���G�x�<Y��1�|z5D�5"��#EGx�<9�'�Yh�ȫЫ��k��ɣa�y�<	�o��y�CA�_����L�q�<��eODhl��3	��B%8u!Bq�<��g]�S��0�	�<&0x{�G�<�u�\�u$�B��J�B�:=��^G�<��O>ܺ������	RƝ��!�A�<o@�k���f�UM�<�S�<Y�ኙ
�-�u�X�|�r�����Z�<�Td�/C��! d��/�d<�p�EW�<	��_�7��X�h <u$f�	U�U�<��L��`��t/F�df���7%�k�<!� ��,ಕ��%��D���A��r�<1�,�K��� bA�a�ębw�l�<��c�d�[���n�\@B0B�r�<��Պfl��	g�]�Y|��
f�<�&�D�0s����F��oJ�u�'�b�<9cH!dչ��ы7Δ�k��E�<�C�G��PHu�H�a��I�<�G
�3x/�q�	7 $��b�B�I�<�" �rE��:͝�/�!"�E�D�<1�h׼j]9D�?�� }�<���
� ���P"j�9���B�<�q�@r���+L�-�܉iF�Y�<)���X	��m�$���1�+ZR�<�PC�&`[���M#h@��Q�<	�l	�b]�D��Ls��RO�<��
C �89�G�:�hE�<�bK&[j�I�۲8����}�<�n+nxޕ���_/4B�l�|�<���Fn�S�)�,�R$�x�<�F2v�u#�X9h�\��fF�m�<1bN� �줒q/�<!@�A`��c�<9�(�
zl{��P9Z��T�I�<���מ`�\��F�A!N��uC�mO�<���!iٴ�p�A(���B���C�<!��"!��I7A� �:Q:���G�<�#"�<UԼꅎÐ�豔dC�<�C1,x�BU�6�thWe�{�<頃 �4XQm�=DR5��z�<� �W���"�ΥKi��!gD�P�<yJ�9=e�� &�Q�6$f��7!D�I@��,1���hR�B�t�j	) �>D�,pAa�t1��TK� �hU��=D�H��"h~�b�$G#-�8u;��=D����U�]�ap��0#�&�'�;D���V�����p���� ٫78D�����W<.g�)S�)\GR���&7D�`Z�	���fM�� ۲�u�	0D���#U]�"%�Q`�0���o.D���F�X(E�$���"�m��ka2D�(y�d�;��m;to[�e��@G%D�DC�ő�]l x��^��R )D���b��eR����˜R[�$
��$D�D!��'�rH��ȇ�&��PrԎ/D�"���NQ��K�d�*��"D�� ��D�ʕ	3Z�� ��k#�� "O|=�c��53��(C�]����#c"Oʁ"'���eS��൩�O����"OZ@�l %������]K�e@`"O�m��B����r���
&h�"O����ȕ�;����o��.���"O��$�j�~�AH[�[��dX�"OhÄ�.�*0Rq!I(Č)ӡ"O�|(A�V.LZPY��	.S�!�"O�D�� $�a8���!�9�"O�Q��N�5^r!4��� �0X@"O�5
ƪ5��8HX�$�N�b"O���ц�(UFI�GS�P����p"O�]���M�\� 4����2���"O搘rA�5%H�&�у���*t"OQ��BQ .!`��� Y�X��CG"OVh+ANp���ʓ1l�%��"Odܸ��&9c�!���ڀRH)p"O�i��� a7���`���M= ��v"O
����;*´�WN]�g74���"O ��L�;C���MA�X.�ش"OĘ���P?Ct0`�,? 6��"O|Q�B��9�<����*G ���"O�%��F�!�vը�D:@���"O����VID"H�j��L���!"Ov9	��[�w�~�w*�+��䊅"Ox���ճ[�j��B*ֵ$|�)C"O�2�EĈ������^f�pJ�"Ohe�Pk

H�f1����=\aN�t"O��-'8Br5��C�v�6�"O(d�wb^3Uj6y�V)����"O��k�(֟)P�"p��h	@W"O�-��EX�xn|�uoݹa�(�"O�X�v%�l�X:2�X�YZ�C"O�pt��/��M�	׏}v���S"O@��sɝ�	�@D�4��we�]�q"O�cD��t8�m�C'֋2^�Q�"ON,��@,ws.�@	�#fV�X��"OD9�@ ٓ/r|!�a�q8R�4"O
��K@
	�V��2��$"�y��"O�t9`鍻vg�A;���>��0"O4Q���4.D���܄L���"O�=ktژC��Р��)9@���"ON ������Bb��"EG0�
�"OġAa�
7$`pM*��E�@�q%"O6�H$��6Y���!HV��1+C"O�D�+f�C��!p}�|ce"O~�ca�؁[�>U��
�Uon$,�yRA��bXi@D\bL�$ʉ�y���$�X�Fd�[�>��2bZ��yb��,�gB�5V&��*"���yBi�����UdXe�%r�'߇�y�� �� ���I�ک� ,Ʈ�y���*}Ϝ�R�ȏT6��&�Q��y"k�D`��j�F��A�`˗�y"U����K��9N,:�	!�y��ڴnxF�j��6�����y���(r�d�2�A7���U��y���&�0<�j�4��]:Վ�'�yҌ;,`T�&H�&}�����ء�y��[�O��a�AR4XH̑�B��y��;p���	��ј[ޚH`Iҝ�yb�
]�VF�[���R d��y�/���\�A�Ou����R�y
� ��"$�NV�����u=M�u"O��ٰ@j��$�EJ�3\Jɩ�"O�x�$���/Pr@�wh�tOV� �"O�P��%/!�DY��C�fC�]�Q"O����.�%:�.	��΍k*�U�T"O �4��.{؍�̖~(���u"ON=���MY��D�6��`�Ш��"On��qk(`�������OEXAxd"Op8J�)|�(����;>�+�"O(5�0���hq�䙄U:��:�"OHA���)���hve[$h`x"O��HE��^�X�j�;q�����"O���n�y$iB�	ʬ�V�p�"O�ųÁ�Y ��
��^�1���!"O�(��ߦ%���sg�$4x��R�"O�)J�kG"	�P��A5Z�h��"O�Y���)��ɛ0��_Rl1�"OV�#���:���%E\BݼD��"O���%-ߓ�h��J;*���$"O2��#㜜fhe�C	�1B��)�"O.��2��z\D�UG�b'�Ȫ�"O`��3L�+O� pL^h7����"O��pd�޵)��U��K*@��0"OF����K#o�ZL�sŇ= Y.���"O�бp�a�b�A��D�.Sh�b"O�АT���`����/{q�P�"OF(IPm��:����BO-sL`��"O�xP�΂�d��f��U�) W"O�be)<��!:�$R�J�!9u"O�����?Ih�@�CZ?S@D�k2"OL�v��!r>�ц`ȁ�~�s�"Od!
�O::�#�/�(Ōi��"O&Q{3.[1���X��U	,�� �"O��$"�|"~i��צ$�r�h!"O H!��V� ����,z�2UC�"O�hׇ֠i���t�[lp�'"O��X��π[\�=�6@l	aahL*�y2�WH6:5��B1|�Q ��ybD3C/u�0��u���#m?�yR�Z�d��E���W�l������yB%D%4;���_/v���Ö�y�V������lH?O1<q(� (�y� �/ ݮ���䚬J� ���<�y��^� 	�D�v/>>l�X�#�J��yB� ]מ��\Es����*	�C䉺Zf�uRR�X%|�х-K!
�C�ɵ4N�PtM2<��XSA��D��B�ɲ7O|�JA�׮��f�k�B�I3*�T E͘M�0!���3N~B��&r�h]�!��zchx���gFB�	 3�� 9��*2��x!�A�W�
B�'D��m��o�uf��(C�.�0C�	�M����Q��Ee�R�K	{C�IhH|�����՘�F�m
�B�ɾAd��O�V�DY�X&�I��'	����Rwv-�$|�j��'k�<xS2;ıc��΅r��i+�'g<���L�4ܝ�!b �3Y#�'��R�T:�(B�N%/qV|R�'�Y*3�	�|V��P�P()����?9X�$��a�p�0H�~/�D��]��	�5 V$z��x���T�N�z���M�ؤbDBB�RX��Z���� D'D��t���0�p��a�RD�#	$D�� ���hT.#�(�H�I�h�Bp"O8	r�KԧN϶����%R����@"O�q�'�mu%��$Q�KG"O�И j��	����Bպ8ڜ��t"O�aP�!D/,�`MI���.���"O18�-N�x����D�O���"OB�I7���tД�0v+�3:Px'"Od|�Du�2��������"O\�5�]R�2l�@�_�ʨё"O��t���wp�޹N�>�� "O*Ecy#h�S�
\}�Е��"O���g�7�
�[@��m�.�0�"O��
�@����@AA�q��m�r"O��B���b���aϪ��$Ѳ"O��*��Q"7)H�C�ԝyp�y�"O(�����&wtؖ*|I2F"O�tR�+SYU�����!���4"O��iv�PT�>�I"g�#��)�"OT����Ne���r� P��Mh"O~tAf�'&�������>���S"OJ��a��)�Pڴ�I�pvY4"O����d�x���T� 7L�4"O���2CJ�K�6��(�+&��ʐ"O�z���$#���WɅ	#j��3"OZQ�t"�&O@|���]:Ωxp"O�)��y�@z�J��Vﶭ��"O�$�@��?EٺB#������W"OĐb�#�#y���s��'tR�"ORUsR[�#�v嘖�A�&���z�"O�h� ��u���R�Bi��:�"O���A���?��ŒK]� `"O0���(&����'���L܍s�"O�8 
�Y��l�,2`
(E"Of��P萴AF�ܳ����]�Ę�"Ol�R�ޒT�@�h�6����T"O �y&�?��b�س`m\�j"O���4��0!��H��ڵ_�,��"O���b�Q��q�w�:'dz���"OrQ3��$���kؓS=�\��"O4$jPFY�JQ5;���X���%"O᩷��B׸dAa�X�s8���u"OA�W@�t �|#%o636�:�"O���$j���x]�Tn�+'x�Z�"O@L�eJ4pTXҡ�&}�4��v"OV���5#-��cԗ..�-�"Oʽ��/�d�l����D�eXLj�"ONEs3��ePl�jg�۪�����"O�x��Q�S�a;�C��P�ⱃ"O.���V�:��d`\L&����"O4HXsl�+!U>q�r���5�.7"O�8���O"N��EJ�->T]�R"O�̻!��W�b�Ƞ��?#�!j�"O��	����4�@�	�%��"O,i��F"�|���O�x�#�"Ob	XF��9R���`H�S�"O|��� ݧ
7�����ٓO=���"O�Y)�ύ�-�(kGd���<�C"O��H���<$j�ī�עf�3�"O.��p�C%\�RDB����XV"�{�"O��a�����Br�Ğ3�.�+"O%�#�+s�0���R�Hmٔ"O�A�FӪc�ƭا.H�!��e�5"O��woA�n���#I��N��1"O �I��ׇ}[� S%�ԚOu���"O� <���QLW�|8��+a��|@f"O�Bt���k:��JJgʠ"O�q0��.� ȩ�H�.s�r��$"O��e�	 D5ܤZ���5:��G"O�I�&gP`�$�7.Y%Kz <��"OrMa����s�Z<E&˪Xju��"O����h���$�^�=gΩ	�"O�@���@�,iI�G�לi)���"Or�{ +�4Q����R��ѹF"Oj�+p&�5xPީx.,`�B=(�"O��j�M�h4 ��
A�Jz�1"O�!	ff�
&���ٱ��t�Ф��"O4�;��׆���B3����p"OΉk1m^[�}��O/�$�F"OִQ��W���q��ʝqu��2"O.q)P/ ^J��w�ʧ3YB�#�"O�I�V%�<G�Њ�-@
�F݂�"Of8#�IO�fLse�J�Vq�� �"O�͢��ǙIŊ��g���2}�$""O�ɛs��L��Eys�H�pg����"O|[%LϫH�d=S�Ƈ7�|�&"O���A��J��D������ �"O��6�J�y��p�gÎԠ4g"O��j K�3�j����;m��;7"O`��`���$�R}8�+U�T��0"O"m1�l@5k2�Yh���V �"O~��f������æ�ȴ��"O����ҙX��  �v�D"O� �q��Be0i�oT\�ݸD"OfpA#�|�J=R��A�YV !Y"O�j���>)���(�.+U�Z�"O��J"6Z�|����Ie����"O��D��ug�%z�M�>�Vy��"O5ȁ�+a� xs._��jIۢ"Ob�8�R�ВA�핡(},t[�"O<(�K!����TM�1N	*�"OJm �`�"i��ܫ�I�#�f��"O41:֊��'oD����?�z���"Oh��"��C�R��N�q�"Ox-�!Fb�m���Pf��t@\�<q�!�\o)���-��
dGM}�<��"���R� Í-F�*".`�<�	�?��jD�b�rl��w�<��P��l�pJF"@�jɡ��QH�<)�Jď�HE�я	�sr��P��[�<��m��q.�0/	�1 !XS�<94�ėn>4<k��V'�1�B�v�<a4� �nϼ�yШN	j�.��N�w�<�g�ئXDҰ"󇏐)�|�5a[�<q`\�@�D�*�c�5'3���!�U�<�!,|n���
��on��c��Q�<q$�v���ڃd�
�������X�<����-�u�BH�t]�El�<a�c�"݋#��T��jS
�l�<�֦�Z�`�����W�D ��DPi�<����i�b�s�A�N�X�#4"�g�<���s��טB���{#�g�<�� �6B'����V�D����^�<�
LHvhx�V$B3�<���S�<�pi�p ��s��A�7?N�S0��T�<G䌈?��j���C똭���S�<AR��uV0;g,��ZHJF�<qB��r�X����`z�`4bJ�<I�kOl��A6(��c*D@�	\�<� �#6ꆧs@�h��KK�68�a�"Of�ʰ����A� W���X��"O����%	;�y�@�ې�d1�"O"�V�� ��M)C���S�j��"O"�JW�����4ף4�d`e"O���5�O01b.T��cQ!	�\�W"O�h��*%���ӡW�=Ϟ}k "Op����^(s��˃n�Gi
�R"O��vK�?}�p��L�0cF	�F"O�0��ك/��Mj����Kc� a�"O^�h����=l4Wa/4Ot��2"O�P���g�Ȫ��֠79ft�"Oz-��J��G�r5-�>	|��"O���B��8۴e[�̞Q��1`v"O��B��LȌA�	��T��y��"O��z�c�E-<l)t��B�$�"O�͛=_a�9�rk�Hr$��"O�u��H
<V*�[!*ɜ1Vs7"OF�ŊTx�������-�ڄy�'��$���A85��{2�H�x�pz�'odE��gGT�r�H���m!X��'�h�{�
�;D�	�1AJ/i ��'ID��s�@-V���`�<6϶�X�'pް b ��vڒ\�g�_�
��'���b��2$u���엟M���
�'�bX�._;6DгvbޘO�<��
�'������)B|+G� @�BLy
�'�� !��
,�F�Z*�
�2
�'q��:���\e��	�"�$p`
�' �5�7�:/-��eݫc|�ո	�'�V�×-�$����;���KK�<�Ui�?5@�!��8�|�2'�H�<ɲ���D�����R�B�C�E�<A@��2.���B�yI����i�\�<��E_Ba1E�/SST��V�<Q�� ���XǯBT?l�zE�WO�<��T�&ք|��
�m� T���J�<��8I!ܵ�a��/K5
��Z]�<��@)g��q���V?Dd��S`Y�<YEb��i�P��geޑJq4����EW�<Y�b�$_L �Юǲ.�� #��}�<9d�D51�,q@m
.o 9D��x�<y��ޣS�FE;��|z�q�GI�<Q�C�.Р���Q�q�E+�E�<ѳ�_:h�����"7h8*�%�w�<�1g̝~qh��f^� ���9W� p�<�gO9V���b���*������w�<�֯م7�B�s1�õr��M!գ�z�<1�M��<%�AbX5zN
A	��v�<�7��;^��c���5P���r�<�c�\/g�@𷁃�J�NQ0��r�<�����CIP�@)=�4�Cm�<I�+$�\q�����E�6�K�-�R�<�TQʜY�̟.7U-)CAj�<�!�
d�,�څlϓnX�� ��Ai�<Y獃[�m0p/˫}/p�Q�_g�<����:`E܌���+T� Ҏ^g�<��g�5;��aF��jC��\�<�fLC�������aܸ��@Q�<d]=�|�c��w�1SeGM�<�&eЉI9�|r2�M<7;���!JT@�<��D�c��U�^��ԦGy�<����qxV�2rJ�c��I�<ip��u���x�R9���7��A�<� F��F���+�lP0��;	�h��"O��j�n�
��# h��s���@A"O�@�$�yI���bGGe�L��"ON�`���0@�[�ݹL���"O���TE�T0pf_e2h��"O��v�5Ovp��E�!W {�"OZو.ںm���:�Jŀh�j�R�"O��IG���`z��aD	��E��h�A"OB�@ׁJ�m�4�K ��
�Li�"O�k`n�S,TiS���4*_P��#"O�	B�D�dF��CO
����"�"O9P�dКw��Iюݱ�"O�H�WHŸ�DJ�+Ѝ"P
���"O~p��cݴ f��34���δ�"O��A���
Fe�d3�\�Bh�iC�"O^!����"L�S��.=n�sW"O�%�䈖�-� ����@�6"OD��%ĝs֨��Զ��8"Oer@�2w���G �Ҷ0 �"O�Ꮡ�H.A��i[�h���ۥ"O����l^'P��˗�� eo�l�"O�0���`����oW\P`A�"ON��l!\�L1��L	:�y(6"Om(���b?�!V�Ѝ,$y�"OP�Rr���5g �"�DZ�R�2b"Oj��!��
Y�+T�ٗ2��k4"O����X�{d�+#�׍]���;u"O\���σ$I ��i֊�1�~܊�"O J��G�Sh�!����&�t�I�"O(A��$8�!�0�G$�(ݚB"Oh����CDy8��0k��R�"O84�D��$��ҡ�6��X��"O���k7^�2xJǠJ�iu����"Or�R���4#��\sq�~�5Ns!�d-��%�0	��{��|�dB?!� �	ǃ.[�\��R�X;%�!�d�-p���*�	C��@2��?c!���>iij��$l� Ka!��7(�j��vfĿS�ν�4 $?!��n첉�拟�nh9�h��!�D�m6X�U�BV�V]���غ�!�uƾ��+�sb� ����!�
�mh�թ�e� Q��A�f͖Y�!�$
��ȋ'͂$��T�&@�,0�!�D�#E�Y�$���\��e�#�͕P�!���r��ߤ6l��	u�Ϙe�!�^2-��@�!+�IW�	S�O��q !�d�Q�d|���?��5�^�!C!��ߝ�>�*Ӭ���2ДmҘ>,!򄌑5+V@��D�U;<8Ы\��!���*��qb�,99�����T"O!��V��}c ͝M!&��iMm9!��u��E;v�2`�{��Ơs
!�dK>\���C �N�g���CJ� �!�94V���%RL���B�D!��)$�B����!bA�t#���0e%!��P!%����&�&FE� r�&�!�D_4�l�j8��M`F�Ҧ�!�dH�W"�(���W9�Z3��N�"�!�$�!D, 2lKqP@X��\T�!��̽i�i�B,Im�@�,F
um!�����NF�,iJ��B,J4�!�d�
4��1�����Z	�R�Z�j!����̝�qF�<[S�	�BON�\�!�� ��N��M�;â��Tu�'"O~���'�8	����BY,��"O�mA JK��&�#����V�f�Q�"O�	vOE�Xe��1;ך�)�"OJ�
�`P����	�3�:)��"O�ٓ���PAj�ruI}�\4��"O��k��\�1�������%�t"Ob�U�S~���W �h�����"O��PfbK/8�x�%��9����"O�S��8���ć+���p"O�cl2'�Ո�ܪ^�`��"OZ����Z`�ҤK�{~r�
F"OT�#��D5ot\أ��5N��p�"O.�@$��1�pݰp&�6C%�r�"Oj)�jJ-��iJ��жb
��R"O^1P�Q�	!,c�&�I ��9#"OĨB��S�tL�$��-�Ҥ)�"Otu��ژ�BP ���0b���xA"O���@&�f�*Ah"+Ґ{�V`��"O�)R�A�NK�]Z�i/U�8�"O2�cw�P�gb�rfi	"T:��u"O:��� 
:�`�Ҡ%S?WM���"OVEz�a^s�����)�"UK�"Oꬃra0iq����M�T��D'"Ov�K��� �r��2��$:�!�W"O���KQ,=��i��]�(9FXJ�"O5a��F�f�>�����;G.�l@3"O4�E�?(N� 
��v��8�"OF�C�!B�K���k��H3�$��"O��L�<�����	$(=F�ط"Oj8�JO4x��F�۶z&0�Ȁ"OmI����Z�^=�RMF�"O��N�2�(�g�ڇ�P�P"O
h�1���b��ۖu�B�c�"OZ4�F�	b�"�*Z(9w4�b"O�u�1�
.��Ui�iW�uJ�:&"O��g���ހ0�ciQ&f�u�5"O�b�To��#��K'��8H�"O��A��8ʄ!*Ë3ꖝ�"Of�F�$��l)D��O��x "O �[U�F�Z���$]�Tz��""O���m�C�D�� �4uŜ4�"Ov�(��8��0���^�:d�'"Oऐe�-��URu&ґx5�2p"O�m����>Aaf�2P���q"O�.ќ[�F���"z��3�"O�"v�eW�����>5"��"O��zǅ$1Fh��A�y�N��v"OL�^�3�8�1d�F�\����"O���L�dxST�>h��i�"O��	A��+��%��
ܾq����w"O���$��)�jk�'[��<Ba"Od�E��=x�|�&H�/i�J�c"Oִ���TYqF\�F��X�"O�Q��Z^~���Y�V�l)Q"O�$
���,|0���E�UP�"Or@01����S���Xi��r�"O�H�e��R�HųcD�kkd��"Of����@�Ru�X*��ҩ}a0�"O@�q�
��_����h���`�"O&����3i	�A)�!����C"OTe�5	�6�<��&ҫ=�
嫕"O�4��K�.��&��q��5��"O����P���L�E� ��=�#"O� NE�&�΁7R0�q��?�b�hF"O�@�e�:��!���g�~�"Oj�w��+9��%���	�Х��"O0����	�%�"(8�NE�]ͦ�:�"O<ܺ�̅�8��]	R.Y0��*&"O�$�eO�Z&y��.��YW�q��"O���Z�~t������[��bq"O�[�*&$�~��A�A2ap"Oh� ��?h{D`�nY��ؐ��"OX�.':��`�.6�lD�E"O\��AK(�$*�fɧ<��R�"Otɣ�e�[p<����ͺ��"Otw���!Ȗ�Kq�(v� ���"O:���\�825 vLy�Z��"OV�2$-P�A����]+l@�cW"O ��fj�0���VH�n��`�"Oƌ����Sm�9��Y�y�Q#�"O��
ޠL��(�J/+gxi��"O�)*"(
�B�$���f՞���q"ORyxG��,P�8�)�˖�>;""O����`��s���ӫΤȀ��"O���'^0l $�R됿oJ�r"OȨh�	�0tHI)p��(4!l��"O�	�I��R�� ��y���"O��g���C{�X:qJ�x�$T�@"O,� �U�ndsvh0`���B"O��+VC� ���� �@��,�s�"O\$�E��R�<�G�=L�u��"OԃbM�	�D��&^2�$Q"OT,�A��E�t�dW�r
jii�"O�mY��۩dn�ʆ%�	T�\Y�"O� �	�e���Iwf4��P�r"OH-8�AV<V�@3�ͽ,�z* "O갈�����̫R
��/߄�q�"O��c�K�j ��W�
�p}��"O\�bLC&\����U`s�q�w"O�)�Rߺ�{��Qe�\��"O2]��$Q�f���̮����"O��U�>�  ����B���"O�1,�oΡ�"EN8B��
d"O��$�U�]�1r��gZ�7"O.}�qHT;zG<l �T�=`�H�F"OB����c2 %��$ѴzN��"O����I^�*ԠI�&��Aت��q"O��ె��G�H�`��F'^����"O6ĂF��6�в�l[���8
&"O|yZ`ꏱ=��Q�k�,�\�`�"OT!��oܦ>�H���\�8��d"O��B�i&zq�E P�jĠd"OVl��
Ͽ(h�Y7בW�Q6"O�yR�M
��Ї�D�bgl��"O�PC���+(�Z��E!fd��v"OT�ڕiC� ��y+� ��z&|x"O �I�Ĕ�<��K`S	
y��"O`�2�瞽PUԭO���*�Ѧ"O\)���ڮ;o�	�%D��0�e"Ox�J�.�yKFc7|�x% �"O��t㙀xw>AZ��[\I���"OFHH�� :>*)�����HB쵑G"O�9"�G�������%!6bEB�"O�0��@X!,y�ۇF۟kSF���"O.O(t "D���#8(l�p"Oڽ(SH����y�zXE�"Ob8��Es}��c��^�v����&"O� �-���\�#rp9��xh
��6"O�4����)~n`��p�:q��UT"O6,p��<m`a3/�D�P⦀��6��#�'0FH(�a�fecw����(9
�'U2@�u�1H�N�*�n^	Y5�8	�'�0���˒�V�,R��%�X���'���r��F�{�$�6 ��c!Ɣ:�'�|�Rd��u&�ʰe� �'����c	�}�*�[�*�Yu~X��'������@� 4�m �O{�|�'j�;f�K�q�2%Ac/�*�N��'�<)Q$�SS��,(�"�	�f$�'!��B�<	��c#Ǌ����	�'J�����6�$P	� �^���'�>�J�(ûm��H�E���d��
�'��M���XWBp	a�	�Zo�
�'��P�	��L� ��^b��j�'ؖ�y&�':���С�J=�')d���Dխ[��%��V�|A��'�Tp��풉[0bl��E�~�c�'Զ�3IC��*����:h#�a;�'���ޛ?��4��e��g��c�'�����M��qr���Mڿg�U��'�f�a�j-J?~��'���M�z��'٪� Θ�:��	1�K��;��$k�'݆���hÛw��X!4b;�D@M>)$"�;�@�<�}Z�`�5DJ�Z�-H6g����ǌ�e�<��&�";����QCM
?���PM�:kT%&�T�!��������)�g��!�a���8�H���y���Br�O�	x�+&�Úx��"��/'������x����JּY�Z��oAy��1��.O���
��|��;��h}�(˒r�(��M-%�A��'���y���:1�8��	${<�Fm]���$T&"v�̹��Z�qښ���S�� �`E�N��<dJb��"�@B��.6���r	V�}�@�oIi�F�2�ϯ(���̴S��l�%����-Lw��:�O,kWRpq�T�:�}b�Խ8����GJ(��3����	��Q���.G\��P��W�y��x>��J5*�K8�Lz2ORy�uEz���<ot�*��@�P8	��j��>��	O�o������-�l�#��RF!��.0�����]<�����{ܘ��@C�?j4��ա*86���M�/�H�׍�R�4�k����t��G8�y��2xz�0�2����|A5f�D����狂/��C���Ph�L0�Ox� Dy���F�����HF��7�ٖ��=���8x�I�Њ
pd��)A#C��1!#�`P�Z���~�
D��s8��P/�&O��@����<H>�LX��;����]b��H�J��r)B��n���N�?}��iI9:d�����![؀��+6D��9�!L]n��@M���MI�E��?�8��bk̂���JbTVL�3,#�'�y'/K3`^�E
�eчa�B]��C��y�g�,l��|ar��ؼq. h�U]�Xd1�pa�u+f(�����𡰆�a"�j� �
<�zr�G��
X�dÌ ^�Z4JE,�!�c��-br����B�JH����>�<��d�Nyniy�/�a@�(y� �"�qO��I�G����H���
z��4{�$��~i��L�e�c��]��`�0�R�S9�H���Pߖ��/�+Q�aK4��q�>Hj%����܁j���5B:����"�Sj�����LuY�`�T=j�R�m��3�!�Vj}4!V�Ւ.�ɠ���rxq��gS�e�B�@ݏl��eCg�h{:I��H�y�,��#�
dg�ap��Q�z��Y�yʈ�u�$z���cN9E��5�Gj�9X��+#ǄO3��꛲{�����9(P�6���]���TkZ5�qO�]�E�N�^rr����5t��f��Y�����[\��oD:��ڴ���A�ȓ#�l�E"
b:l���o�D8�� 2�G"Z/�x×[��Mq�"��rx��w��<��%����Qc�\�$Kx�	�'	���3�]#4�\�C2���+�ʨ9��<�9��P�D'��W�[hc؄K�G��hOr!�̑�Z�8��xQ�ɛ��'`|�p�
�z���z��9� �UZ�J��gCة2��_)?7f�K�LZ���a�'���QC�(a����լ�+dZ.ݩ��,�$9���C���S�,U�������^�d����\�j��ԦW&$ C�	�aD��∕8cpBQKaR84�V��,�P�+6g4?E��'z�)�K�F��t��U ��
�'�����^�	;Ԅ�4Q0���'�ʘ�RX�'����͋^�|��*S�m����)[�q�!��85��Sa���B��ţ'.��7�!�d�����g��5lت)[coD/Vh!�D���`hX���	��h�ᓾ5\!�dT!<�F(3�@ 8��	{��רlI!�xs�谕KO�,�P��f��V�`B��7����D�@a[��(TB䉽H4�P']+P�0�i ˜)XB��-P�4�Cj
�T �f�QP0B�I�M<l�*�ŗ�,��׷rB䉖\��}+�m��AFI��.ɷi4B�	2m�����ПK&`rq
/.�^B�ɿg�|��+.a~��R�IW�'��C�	�9��1೯T=m����W71^�C��|܀4��Մ4ʹ�XbgX&�hC��$/��!���4p��]�&
YqnC��n��j��:q�b	��GR<D�4C�ɍ�\B�D�0,����KE�t�,C��"5�-��E�(&�@��;l�C�I�*��aG�P�E���Yr��!M�B��3A��Q�H�!)������Ɍ<��B�I�|��BVoޥ�M �Α�k�]�ȓ
Y��AE�K�"��',���FQ�+�k�b�b��@ߨz~�ȓ$���R ˈ_ِ��vɤ%�e�ȓ_�\Wa�9�z���G�-8�\��0�V�R�GU�e}�XBv�(Il��	z��tH��T�9*g��^����ȓ<o-�q)��x�Q��#	�`
؆���zv��M���RB���D:r�cN>Y
�b��%�`@;�z�е�HuɆ�	�<��,D���`�>��Y�0@Qo�<�w ԍ.6~�q2�@w������W�'5?%�7�-e����c�;I\��U�'D�<�`V%]��xdꓣ��tz5d�<���eц5:ĥ�5@%�p�Ňċi�B䉭9;(�y����� �C��$��O�����q���f^RU�e`��vY!���.�r'�G��C��<\!�أH
��`�K�-%�Q�b7#!��}��4���E�c vy+�c!�d�hm �'Tl_�(�$��D!��:I0l�ȇ�;ݎ5�(�-�!��ʰ=�L�s���'����E%^�!�V#,F,���X�3�VY���^�!�$D."�iG�1���8�N8Yz!�$�.Uq@���R7�~(���T!���k���Ӓʕ�4���
�@YQ!��yA~ԙ����0�D)FE!�\"*������]�KdpH��R!�O����E�B�7����.#J!�dƿ/겑WmI�%���a2 !�$
eX@5�0ѹ[��%Kt�@ I$!��60IAI-h��	�DL�<'!��q����g�=E�Rqu�0�!�d=[�P9@�R*i�Q$J�6yW!�d�K��YI�G��EF4D���4d!�$�
`>�M:4�7!$�IAƎ@!�� h,��n�� ��i����4��X�"OayҢ�02�� W㐙W�|=3�"O �sff�`�h�8�(��Lpu/��gg�%�=����Ob���5-	dh$쇨S$\�H�"Ob�떉�xҸ}� a�%(^(��-��o��d��[�a|�Ѱn�L%��ݏ�h�b����<����x��Z�]x7� 6w� �a,"8Lp(y���V�!�$�c��;�+�0V̨z�D?3ˉ'a��I� ə|c�q �Q�q&Q>y�	���U�A)� Lb�l�5i(D����74��Ba���U?z0b�e� i+>`s��ެ��"d\zb?OxlANӥ~����.v��:A
O4�8�HV��Rh�q�<�^�[�i�%�n�Aq*��O^ы��9�0=�b�K/���I�`E&LH���SI8�|�ׇ�"	�֏N�O#�����'��1�/͍��@�Џ	�*!��+C����T:0��"ՎۺO��I�uc=�]���TH�)G���貫4�S�P ۧE��*I��-c��B�I�v����ՙ!���1&��&L�8����l�N�1���b��i)R�)��_��/h
diŇ�]��T)2cY*BB���in���T�2KI�>���	]�<�y �D�/���ë�qx��[	@?��q������x��0OX��� ��I���Gl�8��9�4`���JE	`������!
��!��B�ɜC�.�J�f�)L�傠ՠ.I��S�>9�ڨGP����ߧ[��`9����$K �����?o|��ԩ֦�y�aPzN�T�&��b;�YLX���"i8�[��mA���Q^p�|�I>b@X+e����	�2 Qa0GZE<B Ho��1Nզw#�����Q�j಄�Yv�BA*�b�-,���y�|}R�*C"Y�,ѕ���~>r܄�	+�nQ83d� *`����޺^�,�!��[�@�>́VB�'8E���"O�E� ��q����!a�48
}Hd�>)�#¯'n~4��E0kP
�	5�'�`ň'���h�=1�������h�L=y@팋g��SA������)��Ĩ�Af�O�-H���^�g�	�V��7��0Y���w�R ӰB�2�
ś.$͔Q��Ե	H��#�,T��j���:lNY���`� ��p�݈Xt�H�1��g��ĝ�Yw�X�qߍdy	޴n�|\8�&��,AI���4������ �$
/E�`���F�� ��=aRc�}�X5 !�YD���
'u���늆J�����V�,�+"��8��QxU�Ƹ��%j��R<"#qO�}�#q�E�QP�}�,�'�F��ͅ�x����$�.L(t"��F��\�ȓ���@6M�Z�.���/:�����3&Xr �ׄ3��l#��P����E��Y$ԖxH�r� `�^1�ȓW4��feE�:r���q�$��ȓg`�L�D���'|�8��ō1H�\�ȓd!��u(+'I�Y��I�J@%�ȓ|���('@��P�bir��Ŏ(�zm�ȓu�ԋ���3
%��G��|x@h�ȓ �(8Cq�K�"��@H�cJ"dS\��ȓm�@]"%�Z" ���A� O�PFd�ȓ	�*��� O�F ��+U`��؄ȓ��ّ'%�='Z&(�ge
2g� �ȓG8�`���jh�����9k��D��3\z	1T	]=V�t)���"�r0��o�a�f�1
״�x�I�5�I��E�AC��T"x�~��v�K�Fä���Iy<ա7j�~�+�,�Z�"O�Uq���k&pЃ�9P���"O�,;��XjE��O��P��"O��dĊ?�Xy� c��R�"O��y�$#d��́r
*	��2A"O����#��ib��#M�V� B"O�0��l�")a����ԦG�ܰ��"O�h��JX��DP�Ɗo�t��w"O� ��3N�� (B��.��	�3"Ob��!�F���3�$V	q��}��"O��:�HS>Ov���B��6��@{A"O�f�èq*U��"Iab6"O��B��D�e����i,P�I�"O~IqQ)�h�����
r��"O��F��k�!�W�AV#�S�"O��0'�8۞ �U�\c"O��Ɍ�$*"�Ҕ�(t��8e"ObQ�ƀ�0Al,��U��Nm0"O\�9�
�?I�X=p$�<%�,�a�"O�!�BK�< �y����t��w"O�i+�N8v��a��(�+JF���"O�<���>?�$I���ų�8�"O&�+� ��z��J��;F�fȸ!"O�2��E�����IѦ(� P�"O�C+H�]�(�;ʂ,�"OR�p�-y�d񐗍H;x^|Q��"O��14��r�
�sBlL9.2���"O>$J��*Kx&���+B,'�l�U"O��y��l{��4
Cw���6"O�9�#�֛w�M�6-� Fm.C�"Ol�9P��8.� SL	�T�,r"O:e�#n�1y�✋��]�*���"OxA�a�C���
�%��^h�r"O�gF_���w���u"!Pu"O�L��&�7����Q�E:qT��"O�UЁ!�T֮�`��? mJ49�"O��a�/C�7�L�
�� z�J�p"OB�:!��(W�"���Nݣo�iY�|�n]�n�mQ�y���aȚRm@e��Dެ<��0L���y��0�-0��\
0�p�n��4���K<�BO�%m���'����׹ay�9��M
�s�8�	�'��\�e�%��!8Dhϗ4�8P�lS�Y rI`�߂��>�' d�HQ�r�ָ#eFy(��CO�(�JB ��SJ����J)�X�b�w�p�rC��	=�!��ɸC���Z����p���2���s?\B�� �4�8Z�0�M�M�d ��\���rV5.C��>��0;g-H&
r�����t$���!O2r����9����b+��$Ԉ2)D�8 	�.2A�h��N�}�+��LJ��8?.nA��j	$J!�x�� @Ȇ��3b���P��7�<�nIS�ܰfdJ�uI�EFz�MR�pp2ǄI+PaF<k�EK�&���"��\�3v����%�!���8� ��4k�� ��Q�Ƶ�p��S���L�
03� ��0zps�χ��H�'J�:MtȺ�ֱ/�<l�����y""�*p�<�q�f[�!��k�*�e/D�:g(�m�y"b@�>r���!�O�:�EyR̀�^:�����ݜ$���ȥ�@��=A���_� ����Zv��@���e:y�#� P=���	��P0&G8����`�&��2�J�cڞ��T�(���|��8q�# �&+Z�õ@T�=ͦ�>Og���+C�tp�-��RͲu�wl!� �B0t$��#G/0T$`q�E�q�<4+�b	�t��5;��Ôs[p2���kޡ���X ?{�9b䞟7Y�t�&D�LP,�y堈:�\�>s����ǈ�@�ڡ�.K*u���獊=t�֝0un�Gy��͆C�n�S�H�nD�%���>�p=!�*��f�dmV/S�1���#Z4DH1𡕁s@8tb�*��i2�qD�|J��XG���eN*1=z0������'<�YU���B"O��(|L��a��\4��o84d)��ڇZ�122a��Ud$C�ɍ|���!��<n�d	�ʝX1���i��d~��KƉ'����O�~���d�țw���j��ؓR�t���[�l��
�'������I����v���c�P[�)^~
���Lh�Q�!L6s����w!@K�'*�$�RLU���SfHHYZ>Q�ד2ŘZ"�WH[���"��t�-���B�T�ta��%N�t���w\�" S�'�^��ċ��n��0Z.�6�p�؍{�I��x1Xܢ&$X'.P۷�� t�"���ä?Q�Z�Dɻ���?@b��W�4D�� <�yA+Z�6��lB������E(C����3��J$@x�}� kI\�:��2�+pޅ�	D>wh P��eIwni��0D�p��ey<j�!�|�[-�6z_q���#2lp W��q���W�'���a��[�� �W��_�����e�b����Z}�i��M-1���7�/�pd�d�.1k��bP㞌~aa~"nR7}<a%T�59��!�	�	��'�>��\�!h�l�Fʨ'iv4�K?����=*�!a�
X�.]���ybA
�X/jm�iԛ%�ԍ󤃙�$�\��"և3�@�I�O?�IS����/�/�>�	Ƃ�p��B�	2��c�(Z7>t���v�j�I�p�D٪��K��p=��+�.i�x{ DO�#+�]�f��w�<���K���7��0A_� ��&�q�<Qe"��Ri2�y`�C�b^��c-CZ�<Q��P:7H1 #�Χ@�^U�C�Z�<IP�S
|�P80�T432��s�bEP�<IS��7*t� DD@�1��pK�QN�<����&��E����1Y�&i!MON�<���5y���2@\F����Cc�O�<�q��}��g%K�_Ex�F�c�<��ŗ9d�ȅ0�nҸ,$�E�X�<�#�	5�(�	�C�x���L�T�<Y�ˈ�eDP��4R��I�dD�<iV Qq��i��
݈XY��3([�<I 	<#�5:�j�2&,"���@�j�<�7h���x��Z*X˜�)u��e�<���T��l�S��*{�<צ�_�<9B�P�}T4�Z>l�FI�@��c�<�o��%���ЬE�H}��f`�<YG�T�LeV٠���}���g(h�<ٱ�5=�HQW�I�So���S�f�<�Q��U�Y�)P)���F��{�<�#I\v�@�� ğ�6Y��)3GN}�<�/U�:��Y�4�ڹC^ �$z�<����SS����H-ᕉ�c�<��Ju�lm�T� PT���E_�<a�Hӟ@��A�ǁa��83�_Z�<�@͑�ZnI����9��`@P�y�<I�FQ�M�0�K�"��4���	{�<B
T2��3v�M	U-v��� �{�<���@Bq�VH�:.�k7�q�<)a�������#��6�n�{5�WF�<�!\�3�|Pj��0�:�ك�I@�<Y�c�6�� J��_H��Ѷ#�<ybHd�zD���A����+��O]�<���J���v�@1=�R�	�fLZ�<��
6c҆m�OZ�J��0�
T�<q )�!^.�҄̓*k���AV�<�P�O�Q[���#%فl�8�:t�Q�<	BVcp�PU�O�p*j�Z�!�R�<��.I=)��g�?0�NeR��YN�<)��+����@a@�J����v#�c�<�u��>�4���ʁ�`-ji8��NP�<���1!&�k��E3o��ԥ�F�<�3��y�6�q2��5L��)UNG�<a"LֹQr(@��O\��y�MRG�<E�b��@�G�W� �pծk�<�G�	�N<�%BS��yG
�\�<��n�u���� �֌ PѫHf�<�'��uOLE4�C�bRtZ�#�b�<�S�G��6 )�jx}hPX6��A�<)��V�m���Q�
fr�ID#�B�<��D
�(��E[�DK�,�dx���A|�<!6�2n]Y�i�2 ��r�{�<��.ҷ�*��`A.Bդݰ����<� Leꐠ_�`��C��S�����"O�d��_
c)� ��H͌[����"O�dYF�¹.�<�� @�]����A"O�ID �2慲q/�%iw�Ő0"O��kC�p7#C�P�q� )!�Ȓ��6K_5E|��c��H	!�䀲W�´+��O1,�4,�e�!�D��mFT�r�$M܆M@�N[� �!�۴?�i�7�7/@����.!�>l&�X�3@�pg�ݣh!��M9Qf��A�L>��Ԃ4
Ĝ;�!�D�zj��#�nZQ�eɥ鐁;7!��S$LЅK���	��XY&'��f*!�D̙g���Q��
e�X����T�J*!�D^	3�u�R ҙe�f��M<g!���H�NԘ��z�g�&�!�.;�	p��S�D,�I��!��<`��Y2Ʃ�x���:�5	!�d�|�|�!��	)4	��S +�!�F�B�l��cӾ]�P�yS�Ŵo�!�=EĀ�����Xr,\;�lC-D!���:~̠u��-tb�푲aA�!���6�T0�IETv����.�!򤛮fe �4ϛmBE{�5�!�dN�$� ��7�`6�Z�A?>�!�D�ܙ��Ǒq���g�=�!��ɤ$�0����,R,�AB��(=�!�DD1B���� L�4�3kT z!�$������.˧>�3#���1!�Ě�n'�����L3?.Q�1Ɖ4&�!�d�4�%ʳv Kå�y!�E� g�D! �,t(`�J^&i!�䉨I5�``�*çv�"�:�
T�lV!��U��4ѐ-\aX�JgI�(jN!�X�'�e��iܓ?t��.�v-!��L&�t���P:�d�ʑ�عi	!�d�(=f��+�6,����g�D�q�!�$��pb��B̾CZ�`�����3�!�䂖W ��q�H�'�:����'�!�$Ć�x%����b��tsGR58�!�~ lh��Պ[1nih��{!��!Rh�V�֩�&Z'�E�({!���
b0t	���cI��;^�8$S
�'	@���H$4
裠�B�`���Y
�'�������2,�iA�Em��S	�'�yYoW�=ݼ�!��ɞ5P���'-�T2E���1��� O�6D~���'�Ģ.֏yʲ-s��ӊ^\:h��'��r����T�lM�Q��3L�~���'Z6M!����yT �
!�B�(=�'�2d��&E&x�@ ���(,B��
�'Y�MCj.	�CK�/�@y�'��"�dٸ�xh
�Hґ_��R�'E�y�t��W�(�Qɏ�a��t�']����d	o�^Q����(Y����'M�p��� �~� �R��a��'������
?ل{�3YqzE��'���@�&vo��B�C�5mQ8A��'/b-�"��D�1Q�L
�a��Th�'�
e%M8Mo@�Q�GC�	-�K	�'�X�8.H�j <`3�"7&�-k�'��$���&��8����(D�qK
�'-:Q����3���"+Y5t�.j�'�������.Y� 7,X�k�L�*��� �H��+JQ�%!��X�ʀ1�"O��kv�,0
i8�)�n�<k�"O��j��
� ^� ��V�@���ض"O�Щt�"������4�\���"O� �@�.�����	@���d"O� �Aɔ��$=s���>��b"O^���l�B�ZAH����v�H��F"O���e�:1�( z�i<L��0W"O��V�R:�J���)�z��|z�"O���	�'.4�鲇P��d�[3"Oz�i�E�k�h���*��SF�!�D�֛�Pz��,���|��f8Ɇ�z�͍�9����/3 ¤�%���O� æ���I��]��m�3�R$V��m��Q� �����o���S�O�:��g�֨�쵉 �h	 ���~�h�b��c�ҧ�����	�;1��Z�a:Z��	P��^p�Ա*�>�U�EQ)TS �s�C.k�Ԅ�Մ5Z��\�h���sӐ �ܯE^"i��lXP�؀�xR*��a��O��\MBf ��IkHxش��FL�I�X�HRS�#��|Ҍ{�d�J�������3:>(���֬�?��k�����-Y�?1��0��)�%Hŝ���y�(ς+���8}�J�?��S2_�8���9>>�(ѕ��S��p)�U����d�Ob�����|:��?�"�s�A�9���L�%B���V��a��}�]*��:�u���ghG<N,<�;#��$Olrt�G'�
x�t�����?33�M�Զ�0|B�ዞ[���?L
L�;���	 >�\�{Ѵi �m{��)�(�KC�|,�lB�%X�udЕ���>iGsӀ1RW&)a�a����{��d ��ΓLj=h����y2j�|�q��	-�r��|����%��<s�A�*� za����$�4U1 $�>E��
s�՚�	�%P�����H��y"'-y��㟢}ڰ&�-u�&�T.�H.��a&���!���9�S�O!X�Qn��sq(D����g�0a�5&��(�yW�Qr�/��@ua�1M&��>�ulS�����O,��UB�� o&��V' �P:G�xB���O��pMXЧ�/�~��ŏZWV�9[�����'�lI��V�ul��Q��R�r�N�S�'�h�U	ǯ�L1�G�eg�H��'\r �Z����jR?Z�,�	�'x�e�0�� Rh�@r�֝R�Qp�'|����q�bD�V�XQ��'���@�زo@$!d� �b�d��'�8��L�h0Ɉ�)a��H��'Į99��� �>p�p�0 R�H�'Xd
�;�b�`�O[�M��'�C��!G#�ifG�P�~�R�'p���CQd��L�OK�-�'�0 �%��
�ʬ۴�	�F`����'���aQ�J��A�A��nC���'eF���k_�����AG�*P��=��':�P�BD��P��s��|��'����ށ �TY��/��y">���'���Y@ȠM�}�2a�!�DA@�'���s�g0�,�aa܀E �	�'9H F��֢�*d�9����'m�т�����w���GHH��yrJ��5jCʑ6$0��GȊ>�y2�ů	�p(�����E��Y#J���y�b�e}�vk�'0��P�5"�2�y�J�v2\�f��ug�)�����yB�ۨ Q�B\�j��ؐ���yb`�7܉�f� _�b4�e.��y��l���peŮFqJ��j�:�y":E��:$ƏH�X��Z'�y��O�c�`}��OAf(We��y��	"�h]+#䅫ܢ���h�R�<Q�)(i��i��6RL��xCd�<� P��ţJ4n\4�0̢ ���"O�I`�J`���)B|�\�Q�"OV�B��J8P�$=9D@P����"O��r���n�3�!;Y��4"O�\z��ݠ4��1ʐ����`"O������7Fh ��G�M-����"Op�۠�!4��	�F��D����"O��� l2L���CEE'���"Od����C�cv��QN�m=b�" "O�m�&Dq0�%�D(��+��IB"Od|�p�3;q,X�X

$�R�"OxA�+��F���k��(��ȁ"O��#�ˊ�`����!!�h��"O���Q��{k��ے�x��i+"O�ٕ!λ`�2 ȗq�@ErC"O�H�7(5Zܘ�%�	���q0"O&�bUhH��tx3�@}9�HK"O|c�h���ʓB�7'���r"O�y�#`�3,e�Q��Q�"$IG"O����o�w{ZP��Z�Vl��"Ol1�d,�
�8b�P<�Н��"Ob�r��
�Q	���p�xI��"O���5���J �	ڷgژ]v*��v"OqB�M�)c�C0^��� D"OZ���,�?Y��uG�ƻHj^|�6"O`�ӎB�Z!T	���\;I���C "O��]3tgŔ"#��v"OĜ�W��~�Z0L�-7}�q�"O����4i���O�p9�4"O☈�`��0n��H�L��ܒ�"O&�A��{�d��v��r	:��"O����mҩF��!Ʃ�4,��I�6"O�<A���CH����ovrp��"O&�34g\�Z�pLZtiI� ���3B"O�=
 H\�m�Z�:Ӈ0i�4�#e"O���QeP5d��%HV�ԅ��d�e"Oh�.ϭ�r��T��*�,x��"OPQ���	�t�0��K)Uu0���"OHp�ug";�-����,��q�"O��c"�("=P| �
��p�"Oؽ�ƨ%4�]���^�K�R��"O���(P���T:gL�"O��#�3/Ȥ���@O'L�~�BB"O�a�ۃ�N��쓛H���"O����b�<E� ���``�"O<<�cO� @z��kcK�-k�H�p"O�J2��$�X�9B��1�A�"Oް±L�&p1���:0z](�"O X3ƌ�:��`Е�֝(1 !�"O���Ճ@z*�����f'Z-X�"O,���Eq�<��ɼ(�a�"O�{�eB�o_�����T�=t>�"OցA��0%���1Ѳ�2E"OLhH�o�|w�h�d�����"O��1풠9���������cT"O��zS��y��X��N]�Z~�k�"O*M*ϑ�ۚ�;dLZÒ`�"O];d�A�C��1�.[�)�5"Ot(�&
��{F�
b��Yɗ"OVE8b�S�[$=�bJ��2z ��"O���u�F�]Q�����B�ys&= �"O 0�/���t������P*WHB�I�c5#u�R�c� 1pa�L�{��C�	�(9J�+=B��ce :b(�B�)� (��3�Ӵ	$H����"Oވ�t�&*�q���,B~��W"O�T[ oڼ"I���GIG3�u
�"O�4Z��`Ȩ�[�癅c Tӣ"O^Mi�Ǘ�)� �+�&4>����@"O�\�Q��9E��=#�`��|ר��Q"OiBaO�nߞ$yfo�������"O���\?<'�i2�hߕ
�L�Cu"O��+Y���QM�~�<r�"O��0EҖ4�",����1}���7"O�0�!�qt��a�&^���"O6u�sO�

��u�ޔJ�1R�"OPMx�-K�(3�ř� �]��iCf"O��s$��Z�ȝ�f��g.��"O���ùV�T�IԌ �I�87"O���q(�#	1p`�u钃=:���0"Op��+��QR�8��A�B)��Zf"O��CҨ�g���D2P�I0"OBAs"G�]oHU��-�%
��p�"O�|��⟉9�u��
Ƈ7�XA�B"O|�xe�ϖ(��
�c�ar�"O��ZФk�x�� -޴9D"O�yJ��-(7p@��frҙ8B"OB�P2�	�J��1!˶cp|0��"O�}�po I���3-�3^`��y�/�Lf6��Q���3��t����;�yB��FWr�da�8(kR�ju����y��T�@���6$����*�EM��y�K�p��RT��ga��yHӖF����6n-�reP�a��y�$�<��1��=~���A�y��؍\���X��
z���`s�
��y«��(P�U��o|^\�w��y"o�>}�� c#�&`f|P���0�y�BɵOO����ь'?.$K�j�<�yB
�,Ơ8�ݢ �2uM@�y¬S CE���"��Xv�Jt�»�y��Y�.�[�A��
����@LN��yB�R�,J�c߬}�2�R@�?�y�� 3�!�!o��0�#D9�y"BĹ|_�A�"$�4Y�D{����yBBI�-m�eP��'Q2}��.P��y�_�	�k�Fj��& N��y"B(:r�q�D�>f]��)��y�k�&JL��RJ>���c�-��y2&�#�V���C�#J�|�q����y��  0����D����h���yRn�?��!d�*Qj��J�yB�9]~����@5H�T@�Ņ�y2&�&�8��G��B�R5��<�y�%�T�Le��� <��9SA�)�y�!Bu�0�U-�%*�d�i�����yb@�	WC��@Ԣ�(K��BÍ�>�y"D,ir�"E#� ��B�K�y"
|5��)+[�jE�'&��y� �D�X*`�͘=���UG	�y2.D�]����/.e 2�E�H�yZ�X�	�DԞ_8��+ìH/E��y�ȓOߒ��̔7S�8���I�=1���ȓl_��rU+�8!���
d�X�c/V(�ȓT	@Q!S��AN���U	<1A�T�ȓn�m���Jm����q��/����ȓS��w�H":e���D&,�����&����A�W�D�ذ/߽"TBȆ�S�? .�k*(� �S�(ʜx�l;t"OM(:�h�(Q�:.\�x)&"O4��+��0#�D����eM{�<���L���{Fm��}�5�`�~�<y����BM�Tgة=ց@%A�x�<��߭d�������k᎜ꠦ\~�<�P/@\�{A��?��t�s�y�<�1��x�T�8�.6"�0��_y�<�c'7�F����@5{�j��_�<���ɌsB0b#��`Ll)t�E]�<q/Ƭ-�xL�3�UD���8Ѫ�R�<i��%4����"fNhj�����N�<� K�$�H��Fߜr� 7��L�<i`%͕Z� ��ƅ#��|�G��^�<9��
�#ֈ�(���F���E�]�<��!�j��98�%Y�f��%i���^�<Y� �**Y&��5*J�ة��KE�<��	
8]��)b�1�x x5�A�<�Ǡ��-��y �7�p�%��w�<��(Ǆ� ��Ƣ�5"�]u�q�<a$!ܩ΢��4F�pg�H�<��_�DĒL
c�ї1Dd9A`K�<���� Š �"DD��xӒa�`�<�g&�*O�|�dh�p��V[�<)儋_@�y(� C�<�r4��|�<��W,�³Ժ.RP�4�u�<!��+
Fp���R�^U夀q�<1C@��c��U��H´b��]���o�<�fU�Q	d$��f̰&��X�%�`�<���""�Je���,F����D�W�<�g-R�'z�AE��?20^e# J	I�<����Nʦm�6�:IK2M{���l�<i3N�<��)�_�\����u�-T�\뤭֒"�l��0�Z�r��!�%�7D����)�PlD��j��*|x'6D�h�#GF(*�y+�◬3�4�I �)D����P����6�ִwD�{��&D�d�C�K�Rl��EU�f�.m�1�$D�,�`���sߌ���NƤj��g#D�����
1�L�}��у�"D�d��$   �   h   Ĵ���	��Z\KF	�&��(3��H��R�
O�ظ2a$?�K&�P�4V`��ϔu`�P��Lߘz�����E��6��ަ1I�4En���X��'o�����[B��4x��Q���A6�:Z� O:�$��pK\�O��A�%+ 劰�+`�hI1�дf�,��%�Yfy"ɞ"idԳ4�Ԃ��ic�k@E��~�,��!a��.o5�X�Uˈ�g踙�t���)�˓d4B ٲ6^�����ZH~�	D^ĺx�s`t���1(�.~���_��y���mG�|�2$>��
�����!@�)��-^�@x�Cv��k��12"�!ʓ\��O������+B�����N���(�7O^Y@��$ƫ�O�Đ@�ōe���!K�!,
�
E��Z�'^)Gx���^}�dP�nn���Ɖ=���ӣmC���I,��H����"o����N9 �����f@<r�l�'tBDEx����(^6���_80]�� ����Q�8��}�oTJ�'��q�'���0�"W�0Q���-���@+O�]�����=��'���Aƈ�Z���u�ziY�$�d�'���GxR��<� d�?'��3΍C�ޥ��%�	�C`�<B��x��\� i!�)�	8�������~�G�~�'��&��'�^a�F�i��	���Δ�S��M�w�O���2'����֒~"$��6&�n��+_,6 q���G�m�U�ʂʓ�DL�ԩT{�ɻ/���4h7�D]6`�jdCC�
:v�X�Z8K����˷/�'��$�,�1��'K�y��,V!X��;�i8m�X�3Rb�Z�!�ı{� �  ��A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�ou�!Dy�'�:� Ή�B�\O�|�����<a��$�+q��@rsI�E�f�W�]�1O���$���R�W����FޜO��'*(#=�O��)1�h�Z��K�`)����:o�.�<�J����<4���y`���`KR5��O��Dzr��`S��o[X�JC �+�lԛ�#D���5�^;Ki�e:	�L�� 3 �6D��@C�>y��HRc)ȓD�* �$?Oz��L�r�:M�\�H�| ���� d.���'�.���Ǒ����r�Hp*QGz�~RQ$X�E L���   q  d  �  z!  Q*  �4  I@  �K  bW  �b  pn  -z  ��  �  ��  ��  %�  �  ��  ��  G�  ��  ��  H�  ��  ��  �  ��  �  s �  �$ �* I1 �7 3> �D �J Q `W �] d �j xq x W D� �� B� $� �� �� �� 9� Z� ��  `� u�	����ZvIC�'ln\�0BOz+��D�/\�2T����OĴ�^��?Y�+��?�����,+�q2F�ػ
��<��.ߍ"=��Ù�_,���q�B�w�����<z뮘�����	�)��4B��dZ�[޵�A`�'�H����ԗX� d��!T5��|�'c^�g�T�;j��� �'Bݛv//�����9e쳤��m42�ū7ո��4��"����'CDdl�<�4��	П�����I6 ��s2'�7q���t���v@���X����	��M)O��阸4�P}�'�����J�аI�t�5��]�6e��'�"�'��'�B��!�1���E@f^����vG��+8T+FN)�sHў$l�x6tqS��l �"�c�� ���O�#?�b��6��	�vኧg�Vc�����/HR����p��͟���xy"�'&��'��JT��˕`V[.�8Q��x��`Ӓ�n��M3�i��a�Yo��M[�i0��u���y�Aʓ:��1�MY'���?�`��?1��#�?��Ӄr�H4p��f�>	�h�
{f=��T�8Xy��	�0v���d�æ�a�4��O.�Ĺ	��7a%N%��l	�f��x�
i�2�*���)x
,�ҌZ�qoL$!�4S;��2��B+�Mc��iΖ6-��OY�Mc�U$l_0�Qc�N\��1�մT�bA�S��m(ݴ2��vd��M�"ɩ�hW�CHI���P�)?b�P�Y�p9��__�,r	V�5h�Ŋq �$P�7��Ŧ%��4^Ζ鸔]��Բf�˓4�@�.h:B)��<a8���
�V
�mZ(M�<�ڡm�<۠�ɦ�ܑ�E"�O���2�����(�b��7&�*Lj��Ɵ��?���?i��ɽnM��F�PRr@��P���D�S�	ْ�Gf8Ga��'ؚ��P�'i0�Nx�ߴ#1v�(�
A���d͒}� XX�e�^WA��%�(5 ax2��Φ�C}��ql�>QƃLqb=�v���*�@���~��s��Of��$?��B_�ry�=�b*C�H�8 !O���'(ў�>�Z�T���F�>��еkH��b��O��Gש,����&�O8��쀶�'��O*� ����K��S�e��ؑ�,EN��u�Mv�<i�阒fr�ecp��'n��rc�u�<�$b���h�!	8�
���F\�<���}����Cj�2�
�k�@�s�<q�-G����"����d-�,�Ӫ�d�<!B��h}��V�;�T�R3.� �M����?A��?��	���?Y��?������ Y��� ���|�Z4��a�>[���1m̖e	 ���HňI>Hu�,�J�i�9���P=j��+x[D��.���f|!��۾b!^1��� ��,Q�������.��zP"G�*�Ҡg�r�qᎁ	H� e�u@]��&7͏FyRHۮ�?������|"/��(ؐ�u�̌9�(hs��;9�'���'3�������J��I��W6$[4悁l~4������$2�'�����D�|�������H�⧄�9Kn��	�fQ?�I�1����ٮ`��)X��2/Q$��O؏<�!�D��$�ɺ.��#+��9'��8�!�	
<n\x2�ن#~�`�ʈAt!��UT��'���&pB��A�2a!�d��}aF���BDi�+d���E��y� n���'���I�Ib����t$F�"k�0��'(�P��'�r�'� ���BO̓��*4��Nƾb�@���H�I�5␤أ;sax"�H9u*F���j}�2��S.��� $K�v��£=5�F���Ȫ/�џ�ӡ��Oh�o��M��I�(��6m�-6�볅E������?���?i���'��'.f���evr�S�ĴTV�J����>�i�X	���&I p #C�©\�+��d���`�n�K�5�	�?�:�F�4�| �ʀ%&���� �p�<Q�!�(K:����c4�;�i�g�<q�ժy�Nl�7�ь*��z��e�<ل�_(��(�7-�l�H�2�ƖV�<��KD�r#�@AV�'�X����T�<1�@L-��W�RԦ�ӯ���M���?���@}R�Afd^�?1���?�����"Lˁe~V��-R5p���j�\<��<q�ᘛi��N�elJ�+qQ>�B�^�G@Y+fj��\��,qI�8L�(�b\-�yB�	!��1���y"�˳1���r�W��`!��V0�?B_�\x�%�O�I�K|�Iğd�ӟ&@�C��"|ƒ�k2�ܾL氄ȓG����4?��#�(
�(�6ܖ',26��Ц�'����?A�'�>M�k�g��\��Z�A|>=A6�K�hHJI`��'�"�'��Kp�E�I���̧zaS`)ܺL���
P>|Q(�c^t<i���#'���p@,w�88��=eD�p���$���xp�Q*:ODɊc������f�՟H��r�j�xD��*�\i�4 �Rϐч�3�����"���#X	~t0%� ��4��a���0�Q?A��@\����IZ����	��E��%��ϟPpT
����I�|"e�L�p��Y���2u�	�4�� V(a�V�E	 ,b�h�����)�r~���S��y0�sEޤ�M�R�*uR�$ĝi�����,�v`:��"'�9�O�×�'�R���b2
 	.Ѕ9�r`��p ܐ���0>1B� >�@Z�����h[��s������C�\�2i��J�88�vC�|n	��sy¢}28��?Y,�HT:���O�=`rL�>'D���Z�o�$P����O$�d�y6f���5(�l�iq�_�ɔO���fT��@#ߛF�q�������ڨ:��ۘ	V*���ʆ�h�p١D�F%<s�%Ђż4�P��Ě��C`�O0��A��^�O ��a	PG��	g�z}�m�L>I���hO��Z�l	0���4٬�Sl۬]�EB�b�4�m�P�IS��	R�!�/+�`�v˗ TlZ�;�O���O��蒋H�g�$���O���O��nP
�d����!8!Dр��m�*=�P�!<R�oZ8u�YV˘~̧��~� `Ku��.@�T���E?a�pH؄	I/d[����43nd����U��Odl��
��yG�r�UD�"h����i���k��������'�ў����L�eK,�)I!4�ȵ��f�<��T�$f@�"Ăڱe.�0Cea�Yyd/��|2���dL,9�`�; D�7��X:U�V!Q���M�!V
Z�$�O���Olܯ��?a���DhG�.*�A���T)F�P@z���Q.:=�� ��h>�I�Ͽ.}lq��	{�t�R4��9�X� �ƌ!Z\� +ؠr�~Q�Pɇ!ϊ���'��UJg��,C�4�3g�,hljyc!��#�?�i��6�:�I3��OK�AّaM�B�9+�o ��p�	�'�|H	"BB=G�h�k�_	TlթH>�e�i��W�0�P�ތ����O�T��?8g~x�F�7T�B���O<�dCj6�$�O0����Q��.D����@������!�.�%+�M"e���`dbJ���O�rJ�''�X��ť���7-٧at��*��H3H�P� 2�R�`cZ�v�ȰeYj��?!�,Kşh�Ii~r�,[���O�0�
�Qt�J�䓓0>a��T/>-���Q�*�ƈ��OF������Z��F��{V��@I�|����Ify��Ѱ��'��P>�+�Ɏ��D�v)�E-��`��?F2y3�`	��I%Xc.m��",p/��e/��?�O���^1�Bv���}}Cw��zk�O,Q���S�5��,@�㈣}���L	Hnp��IRJ挓sG�d~�!�$�?����h�*�	���"�b�	*�����lkdC�I?tP�M��|� ����ц?�X�?)���3IC<=��H�8`�-��O�#�&9o�矐�	韠!��] ��<��؟0�	ޟT�;	t	qd[>^X�`̓	u6�ӂ_�&+�u����/>8��a[�'%Y�'L�E����VrΩ{�.��c.��ۡ�ڵ�`�)w��!S�B�s$�1��O��O%�̎+�L+�˞� S���B�'_�I�nA��D�O��=Iơޜ+����@�0KT(E2�+�y" �,XY����dF�n�N B7DX#��\l�����'���':�ƠRE�V�k施���6���$Pd��b��hQ�(ẅE�D���C�I-G��)��۔#�bQ�w��uf�C�	�Q�(m���ϛ)9d$PG܃p:�C�I|�D�7 �w�.���[W��B��c��Fe��{���阏[&���G0$���Ք�@�Q���e���pg�?�!�R��`����1Z��`�!��11ʕ�i��q� �{7���U�!�D֮�*�0
�~��4�G��e�!���v��0C��H���@��Vt~!�$H�~����Ԫ1�Ե���"ў�3��-�v��)ғП(͎��% ����I�ȓA[6%��f�{��}�3d���L��ȓGPp���
bI�>{4	��J
\�q���<0��t��$�6m�����	`T�q  ��&P88�H1n�e�ȓ�xjF
;���ps,�n�Z$�Ii��#<E�d�ȓ
-�!�D��~�8pv#Db"!�"|�\x���{�B�Ï��:�!�ę�|��q���U�е2��-5;!�֪9��40�N�7T����D��&�!�J�@�(:3����c#ֻ@X!�Qt��Z�K���ÔC�VG�ɑv���ĈfL�ZdBI{w�)
��~,!�� ��R�D���(;��̫7�y#0"Oļ��ya�P�f�͆�z�se"O\�"�,�<Sz��	\�O@z�"O&��80��EJ�g�jV��@�'�pA�'t
$
V��ED d)֋Ӫt@ �'�B�{�
R�f]:E�A����
�'�-�e��S��"���(:��	�'<И���F�m��	`m��HTp 	�'5B�"2�1h0y��A2n���'o�9�'Z�3��huh�j�����~�Q?	
PM�sD6�@�`�oZl��b�+D��bN%>�.����H��4U;q-'D��ˢ�	� ����AB,�PP�J$D��A��GF���sh=)ԀP�`�5D���Aʜ<_����A$ؚ8�@�F	3D�@��*F6"�^5��Y#c�D�+���O���U�)��RLbr���Ʈ!��NJLR�e�'_F��^P�;�dIll�
�'�p���j�i䱣S�H(
�V K	�'�v�h�gJ�Ew�I3��I�U��1��'�N�x�-ݪ'*���Ɏ�K�X�2�'�R�!�E�^Py�+Ɯ��(�+O�����'b�ŹAkǓ����e�\.�I��'�`�yAjF�:M��职Ѓ^�|� �'�
ea�Ia���i�O~:�'W&��
 �,��tn�B��e��'+���S) �Z�9�m��<�R��
�C�A�*�T̊g��J���S�_h�f���s	v�`�ʴ`P�8@�M��t��+p��P2in)ʄ�	_G�m�T�8D��r�f˸�,\���9�ΑC�4D�`)0c�/b��t!n	�� �4D�L��� l�1D�SI���e�1�8�عD�D�,{l�Ё0�I/%��!�����yEѐG���������w��y�FX�h�b\�R���>`{Wa ��y"��|��cf����]4�Љ�y�$��Zr���%-�'�� �쎺�y��%L�*<�sL�L"���Q(�9�?93BL����0�	�C[�[����c��"32�hS�7D����̀4v�\�ce\���YE7D�Z�l@��|�T�� ���Bg7D���$N�S�h
��Y����E�6D��.Lnd8��ǚ9����k¸R��B��3��ؠ��J8OZ"0��)�NX�ʓT���$N��q�-z� ��sC��p�B� J��%��bH�Cl����ڽV�B�I*4/]q� *Ԍs��T�k��B�	cy���ѭr�fu�^1��B�Y�Ƞ�7��6�d�ӔoQ^������b��d0n� <�aG� ���R`E�<�!��I�h� �˚`w�0�Ad�!�D�&�L+�m�E���F%N��!�\(v�*��u��$6-��n
�!�$Y�1�މ�%@�	h� a���ī-�!�G�!��H�
عU�2�Th^�8�ў�f�7�'6�i�"îGl��3((v����xy I4�VMTM�?Vp��ȓG���c��\�����N��Ʉ�
��h�vC�.��HK@��1dGV���#�>�
�i��e����J�*>p���ȓ.�P���.h�<�c����|���>t�#<E�GL�.t�	�C�~�`��u`�v'!���)B�") �/H("�ܙӗ��X3!�� ���0`�<�&�ӡ���x�z4��"O��S���g*�
C���Y7"O88ʐ�-z�z�*�!Sh�F���"O�@�æ`�F�w�D1g�ȣ�Z���rd!�Oj!u�23Ul�3���G`�F"O�Cd)�su�t�rS�_Z���"O�DH�H��j�1�ÕiFL%� "O�hA�b\Ah���V#[�8:(���"O�$pĨ\6�6�"���&:�����'�HL8�'�n����)|ͮx�1�� ~"2�'�$hv�Ƿx�^�y��|�*t��'@N	X�F���1�@f�j�f�
�'��4���D-2�D�G)�bŌ�Y�'�n�)��@7��`��ոUF�]�
�'9z|PCk	�0�P���'b���ė1a�Q?��1 �/�n� c��	��Hq�'D�t0��n�T�c��TD�`;�()D�d��J�&>*\k��I�U�q�f%D�x�s�O(,N@Ai�ǆ1H)��ZK8D��4�2GWT4�q�}WN�HW�2D�,A�I4�j�s#䈼_���g�O:�Xf�)�'q�ı��	�'aTȀH��3�
�'r�B�/ĨRy\�B��L5/ڮih�'s��1����V�ДM)x�����'�.��`E�@���C=�Xز�'4~l���5g��"��+1����'�N��nH��(BQ�N�(J )X(O��[U�'�4 P��S^�Q+�̷�*]��'	b�tk7��I�\"��1+�'�꼙C����	 c[;����'@,����M8�59`o��	�^ih�'G0�*Pk����X!Ս{���	�n(9��"�x	r�
:Bގ�re`7b�X��p�0��2f�h�f��4�ɸw?���ȓwx,���:(Id�
i�?rb\��b-���f/�n���"���{�ʑ�ȓ$�Z]�Q�͕]���ڥ��B�v�<A@Ȅ&����gE!^q9{�$Xk�'R��Ɏ�I��2�+�P� �"����)Y����ȓ
0T��O_( w���+�'\v�P�ȓ`�t .�'�j�(Jм�@�ȓ)�F��")��;�������X��?~䙂�ݤI��:���B�����u#��e?]n�����8���I�a��#<E���B�L�)s��:&Ԥ���>{�!��i4H�ö"�T�q9����!�Df�u:�-_5�z�Z�Ϯ9!�Dc!t�P��n4P�y�+��G�!��q���cĨ�>h°����Z!�$ػ���SI���d�������'jJ���-=�ؐ��$?���ʕ%���ȓJWt(!b	�@��³/K�`�tA��KA�����#C��:��9<'�ɇȓF���Q���F��]�1\�h�j���W�Ԩ⁮�M�p�!4ok����ɼOF�	��5�m�^��7�[>UI�чȓb�X�Ua5"\��2�ċ�k�nH��A�l��O�3���݌P��u��(�¡'�ì]��U�%�.#�*���o�\YU`�P|��P���z�d���0n̋��)=yT���a��]�AF{���8䨟���1@��bN��#�I-3�lĒ�"Oؕ[��S�YT��r��ϗ��Q�R"O"�@�l՛? vu��ʑ�l�A#f"O� ��2㊕q�Qxg@ٔP"��F"Oj1�a�b����caqtt��"Ol5��܃P�:���i͸�T� G�'2����Ӻq�Z�2�e�b�B��G�G/M/�H������E�ڞ���j�,8j�0��E����a��
Ά�
5/؂l^4��$&��s�3X\���HZ#P�ȓ>�p�1�m� ���S��O �!��q��,'�X	Z�"��HC�7��Q�'ږ4p�y�U@�^�|����u%Io�N���TSz�J���#վ\��$�0ȓ��y:ƭً4N���Үȁ5q\���N� :Cb@+`�^%�@��=�M��z���Ycℕ��@{���:s%�X��	�����d�$%3n	�KZl�YC�@�1��B��"^i�9ڦ�$VD	�1#��hB�	'^���0 N�%W;j0C2��&zB��9\�T�E��&:�(m2�`8L�C�I-��@���1D6X@�K7O��C��+���9s)��-�>�"4ߍ C�=�C*�W�O(�$J�/��	�lqS(K'>56�	�'vf8i�N\,aKґ�5N�6�t��'��T�έ|�h`�Q�P�{���A�'����C�4x�	Q �x�B�P�'i2�* (�O�À`�o<dq�'�#�(�����pX�xu4I��-w�QGx����8EJ��⃛)=�0��qݖfa&B�Lk&��bM��5!�q��Z��DC�	�![j���J���,xV)V��@C�	�=��-�� <v���R��G�ZC�I�C6�]�2)J��z2��6Q�C��?��<S���!]��M*W�]�	�b��IL�$g�"H�F��;Op���'�?�A���F(d����;~��(y��	+�?�t���?a���?�D�x�"�`���L�|�9���yjP�]��9��D�NA���l\i:#>)���,��� �Q­1ˊ�Y�� �zw�Չ��*�J���?hn��W��O��+�Ӭs���s��8X0!C�m*���0?i�iA_?8I�@��z���ӓ�jx�<(,O d{�
S�(�����	M˄E�^�4�d��(������O�]���'��)��e�Q�	�sr���4`&�\�*�J�H$%R�^e�1aUb�i����O�1��1�sFR�<(>EX$�,)�t)t5O��hޟe.�I�@͚)Ph�����Ⱥ[�Ǒ��x�.�s�V>�Q0���-o�f͓=����������'�����v��(T�K�1�ɝ�A�!�����R��B�V*jPPѮ��1Oh����!M�zD��-Rƍ�cK�@��)cF�����[ʐDɱ�~>%�����I�?]�I6y�%q%$Ҥq��$C>�*�d'Չ�M��� �B�0�]����+��C�zh�C���\�|�dl�1P��Q7hJߦ��eb���&�H��

����Z��P�nH,}�v�rC��4$���;?)��֟��	{�'��d&'�� Aw��<����AF0!�D�O�m;Vh�-j�@��@�[jV�2��'z�#=ͧ�?�(O� �jP�V�EyE���#��}9�+�4P�R	�O���O2������O��!;@<�f�ܤ)�Pu�U�K:rؘ%3�f�w�՛#�[<i" R���)��O� KSA�*��BF]6��0�5d�:	2���X��`AO ?��n�����/��8�U�H2$��؈
�h�i�����`E{��
$����f��3>6xZ"@[�MA�B䉱w��cRO���r�)�̆�)p�ʓ.1���'(�I�� m������o>�;ai-�9f�T3(�f��/�O>T)5��Oh�d�O��B"Ύ�e�� X(�<,�)ɠ�u��A<f�2Hc�Y�@܊��׫��Ox�)T��9฻CV�fLs�cغ��%�8X'�����L�?UA�	�M{D��W?A���OX��Q0�y�Եc���s�X�-O����?Z���֧w� �a��}2��<Q�A�1�{QN8z�b-�Q�@y�
�,#���'BrS>QH�@�Ɵ8�I#5��p���&$�Ь�Q9�P��
/d��SF2�pV�I�[X�S֟Nb>�2rǌC�r�(b��Z�^�!7ga��HGJ� Ȕ�DK�DS�tCa�L�u�����%?��Ӏ��c��7�Z.H���aa�4 �'�"����F�S�? l�qȅ�}r�(��� ��b�"O�Y��荩p��l`%�a�c&�I��ȟ5j��ɥx�4��ơܞ�١!�O��d�O�,@���l��$�O���O��	�O�H��5�ѓ�A�&]���Ub�nz���	�>lԣ��@h��g�'��8�&fE$9S��84w�`�-VR���q�V ;!K%���ɂ&^�1B��/Q�����.a�t�\#�<��ǟ8D{�0OB���NE�2(�] ���Qx� �"O�*�G�y���a��t�'�#=�'�?I-O8ԣ&��xR����g�+���IE(T/k{2��e����$�Ob����d�O��S�\T�$�]\���a�0�X*U�M@0�Y(�}��I?c��13��Qf��We�)d����޶F�A��A�LU���	7F��(P�h�A#�"i �5#ˈ�*���ON��Ѩ�<
�&�rF.ؕ"O|M��J���R2@(3�ȼ�Q�q�4�?	/O YX� ��!�	����'D���#��1�(��f��x�p��	".�z]�	�����g�h��r�S��(��7`c�U�v��K�臾w��*�Е�~�0!��r�'n�M�t"C�k��Dۧ;C�eu�}�M�'82ʖA��[n=۔l�		dM�?a���`E��D9��t���E������y���,O!��h� ]��Ǫ���>Y0U�`)b�'y��[
�̲E@�<1��?�K>�O~�=O�=+`��E��� ��g�y*��O�(��K�W��hO:�@�X�vkf!ZQN�3|���d�$o��O��8O|:I\�K%���D�^-�؁e�ѬB��&�'<�̻�;O5���'���O�;OR��ҥD��0���ޚ�b�0�E& 7��O��K�i�O��	"��s��΅d�\c�Bݸ�g&(Ȗ��&�_��d���៴���d��͓�u��'�r�Oc�9O�i�
[�,J2�b F�� }�#��'>^R�'3`����'��Dۍ-����u�a��doH�4gx8�si�Dn�bb�ϟ�rs��O����+*��Os��'����'BzM�G��k8���g��#Em�p� M�O���v�'	���y�R1O��ٗ۟�^wZ ֝)8*���ьY��t��%P���ش�y���,�?A��FX��O�r�'����ۛ+�"�9G�C��ɩ,{g��58Of0t�'�"�~��I�<A�Jpn� H7j=8�)ݯDӺ5�q��{{�i��V��M�'1�u���it�7�A�K�z�̺�����Q`�_M�}�B@��r6
ES4-S.bڛ���5zQ��"h���'��4�'��%\��Ɏ%���o��U8��r�/g�7M��b��'T�	ʟ|�)�>9T�D�����\�z�J����f�<Q�8�,�Ba3n0�\���妕�	Ty�'�.맫��|4d�%�
L�b�ѝ
��PUb�%X����'KQ�d&�b?�Ӡ��~��A�wA�gf��9�4��X��j�'���$E֯y/�ՠ&�	�cD��'� �Pc#d�|���8kXIp�'jF�YG�#k�y򉀻\�D���'V�%�p�`��!j�0!�H��'鶽 5���F����^��j�'8���4��Z��uc�)�9���;�'<����D�/d>�qhZ3����'�)�0���O3��H�K_�uY���'�H|�!�M?�|d�ɖ�f�pи	�'��8HqD�.���HP!�3�t
����Op�$�On��O�3��%l�ٲƧ3���q��1�	����	џ��Iԟ�����|��ݟX��#��>lzfMę�l��U����O<���O��d�O���O(��O\��S�@�6���E�1M�q�� �<[�=nZ����������p��ٟ�����L�ɶU�����D�-���s�!̘b$ ��۴�?����?9��?1��?Q���?��� ��2#�T~ȺF�R�n��Aj��imr�'��'=��'7R�'�2�'w$e��K�1iP@�����s�)k�h���O�d�OH�$�O��d�O~�d�O��#O�3"ϴ�P�J�X�L!�mFզ��ϟ�����IƟ��I��Iߟ<qFb�/�|<[v`�  ����t�7��Or���O��d�OJ��Ob�D�O��D�ofe�F��m'�mцڶa�*�l�֟ �I������şP��ɟL�	�L��I��hɬ��q����/"�Kٴ�?����?9��?!���?1��?Y��q���T��=� ���T�pAV����i���'�B�'m�'a��'���'���&�26�l[�M�W~�y�M�ئ	��ßT��$��ϟ��	ڟ��	��Pօ���J�P �ƥF��U�B, ��M��O���<��ɖ#RC�)���Ȅ#�p!W��=>7mN2��'�tn��<IR��
��q) I�w|VAA�ɖ�� �I�<i�Ol��N]��o�V�	�q��sC�mc��Bׂ��~T�D}�`���t-J�=ͧ�~�	�ڦh3�F/k�H�@
�̟<�'��'V:6M�)��'N� 8MS���l�f@zDY	u��x���t}R�'�R5O�˧P��aؑ�[�~u�E6 &��'�$��F��`p�O�)��?��H|�4��B�
���#�;�$�x�<Q.O&�$9�g?�T�ʌX����R^�(`�#������ܴF��'�7M%�i>����T#Kb�h����gP�9�c�4��֟�I~�t}n�n~�4�������s5fO�/��1p�cJ9��`�%��n�'�W���|2vg��/�RI� �
y�ެ��gy� f�0�{�{2��V�D��q��ץo�F�"��*W��%�'�2�'��d)ҧ{&���AV{9{Յ����P;fq�'&����r�|2V��SƂÍ~���P��C���%JUǟ��Iş�����IKyb�u�Œ���OPd�5*�z�A��°s.�l�T��O�pn�_����-�M�G�i��d�>�b� �]<&? �p�BX�F�tlp��i���h�]�|��;�?)�'�u�H~޹Z�o׻m1��*f��9�V�����Ot���O���O��$�O�"|:w�R�,rA�uO�}|(��ՋR͟��I֟��޴Y��Y���?�a�ie1O�Ͳ	'(Q�d��Z w��}�a>�V��]Aߴ���%A��Mk�'y�U�rA^[��(8P@����G)�/y� ��C?�M<1�Q������4�	ԟ�Р	�0?y\|�'��*���v!�� ��Ky�~�lP���OV���O��	�
�k��֫��Xۖ��1��=�'�~�oc��Hb��1%��O�뷫�3s!n���Ј[L�p�F��8`%�޴]W�ĉn��.�
���#�D\�B��Ch�=@�TT�שQ$2[x���ğ��	˟���j�Fy"�b����cg�5Z��"q璉h������:t����O��lP�O&�I����n�3<<|���Q=::�B�ۦ�z�4K�>��ݴ�~���Zϴ�8�-�?U�Oᠠ2��$N�[ÇY}O�7*V��ڟX���� �	ݟ��j��O^��r�#�C�/H((�Ƈ�;;כV%Zw��'����'��6�m��'�T2E�a§�
#��T�ЦP޴G��'^�OY�!г�i�DG�G�`P��>�(s�*ɝ3����uv���4'��'w�	���I�<�L$b��2U��'"�x}������ߟ|�'�
7PH����O��.$v�[�Wi�Qks��_o���O��o��Mkv�x�+G�P0���� �#Pr�U��>X�t�B5�X�0ת+�)���?�׊c��� �:)K��귮ƫ ��O���O��d�O��}b�'Tb(���IJ��0Q�x^�$��!��D�&%�	�M���O�%�	$p����A�H|PE�'Y�7Vߦ��4m�۴��d� 6�����'"2̀�O7y���.�6`�xUc��)�d�<a���?���?����?!��M:��-"���n��i�������`B�ӟ���$?�	�6-bx�SJB�_���2U�I�/��L�Oz�n��Mx��$`H�+f�|��wC��p�)�c^r��c��B��I�0�	���'�
='� �'κ�7eRe�i�6�]�hr���'5��'z��')�W��9޴*��ER�'L�x9ǒ�q5�u4�	i�����a���dM\}2�~��nZ��?��(U��\�z�HțYo�$����f��l�l~⌇�_���7W��O���G`��x���-gx��#�L�/,��'���'�b�'�"�����6Y�Rw�eQ6nD �,��O���ܦ�D��ğ�����Mӏy���Rr�@`��&�>lÑ����?����?�qC�M3�O��Xe,m��Á?;.�IA�̰@���Aw&�O�+K>q/O���O����Oր�uN&B���	�E��$j�h�OF�$�<��i'��hR�L�	[���]�>�h�&J&X�t��2/̖��d�_}��~�ʰl����S�i�>?7\A�j�h2q��>$�6�3g�>��h&W���ӚK�2��L�IKbZ��7�<��Q�f���P�����ʟ`�	ڟH�	w��OyR�w���eǗ�{��C�A	T<b�ě|z���O^0lE�� ���M�`A%3���_;!���چ��2U���cӀ�1��o�r�4\	�������̟��Pg�V��sbS�ZϞ�[D�'��ɟ�����$�I��<�If�4 ��?2̨�
�8%6R�^*�6`ڧvR�'���D�'��6�t��Ó��� $sa19�r�����q��4ʉ'.�Oo���D�i����T!X���� hhD�r�y@�Ae�Փbװ)�	-+��#��˓�?���9���4OT)�Pd����f�����?9��?�,OFioڿ����I�`��,WY0����c��-a�h<�?�&]�\��Ǧ!{L>��ܾ|4��f��+	� �c��By�Z�K�^uR%[J~*��ƛf*��<a-P�n��A��-��X��/W������T�	ϟ�F��?OB!�V��$*ۦ��A/Q��\ʀ�'J�6m	.|6��$�O�nS���b�N�b`x�q�D�L��5#�*�,�?)4�in�6����I4��զ�'��eh�U�?�1S��&˸4|*(��ҶՀQ�|�X�P���������������q"�SU6P��$Z���d˒��Py�Dc���P�G�O����O����Ĉ�f���;�g�&BT����U%�Z��'�>7�Vꦁ�L<�|�@�~̸;#`ۏ^ �����l#�A�`L�;?6˓6���G��O�|�N>�/O���]�8�!��B�|U�u f��O����OT���Od�d�<��is:P�`�'�� hA�x�\zq� C\h�(��'wT7�#�I����Ǧq�ٴr W�;yBXѱ�S�v]�uP�f�3DԳٴ���͚T���Or�O�� M'�0���īQ�jK�Z�b�'Hr�'��'g�ᓓ&�0A��C��'�B}Z���]�&�d�O�������Ey��~�pc��q0�J�"�	8v�1e60�R�=���Op���O��Q%tӔ�Ӻ�2�30���)�G�8G"�p#�I"N�5;��w~v�O���?i���?��
b� ��G&J�Ɋ� 3�4R���?)(O�o���[������IX�$�Z���$ �'�hXr@���D}��'r�|�O���d��Uk%���r�$2x)@&	E�U����������O�T�J,^5) ��![z�<��n�O4�d�O|���O����˓.���\1s�<Az֌�l�RM�$c؞l4�b7[�h�ݴ��'�R��?�v�Ԯ7�2�ہ��,Oӌu��K�?��"�=��4�yrԟ��{�m���u�*Oژ�B/
j�`��V�E�c� �։�O�ʓ�?y���?����?����� 1���(`�A�F���"X8B\6��0����O��+���O8Ao��<����7}R�[��6�{����|��}��M��1 K��n�Z?a��K��H�� V����m�ɟH�$NK�{b)�L�Qy2�'|�ږ>��#`ĉ��=ž��3�]ş���۟���Qy�g~Ӿ8��O����O�|�'Gӱz�Сr�`�;0�`�<��OZT�'���i���O�� ��=&�le`˰j�&0��]���H?_�@�l���r���I�<��ϓAʰ �&�$��<��矘�	���՟�G�t<O�@ �g��Y��+�� <T��T�'jT6-V;|G��D�Oƭm�X�I����T�\=���C�\Cd��zFd��ɣ�M�U�i�7-�2�6m6?�H����)��b���6�[8e���ۤ�݆u�p��L>�,O:�$�O���қ6�'�2��0ky�an� �NdP��	���?�M+u���?����?qO~�����M�5a���3�N^�u'�J�_�1�4웖�$��'E�����ˢ̌V�I��U�	�B$���(O.m�SM���?�&�+��<��#��Q,��{"�fM���?I���?���?a���ԦY����<����||��3拞�-Ʃ�!j�ğ�@ߴ��'K��$�� f�6`�ɻ|�(9�A�"�e�"��uʘyp�x��� s�-�������AJ~:�w���Q����y���f60���?����?����?I���h�W勞`@��F�	\ΩҐ�'S��'s66��˓?�����GLŀ�����n�p�E0zO��n��MK�'�01�4��āc���cv���j�n
�mJbpIiL8�?���.�Ĭ<����?���?��Z�"���pye�O.RW2t���?�,Oz�m�pQ�I�	埐�	h�$02�&�s�D��(�ctLЕ��HWyB�'��F=��?�`J��%�N�c
h��RV�1t�>D�]�{%f˓�:Pm�O�O>	�g�8g�@:�&�i���N��?A��?!���?�I~"*O^\m��������O]T� �%�h@����������Ms��B�>���iS�|2�Y�1b�3#���x�d��%�j��1o-7�:xm{~��/j��S�x���K��B�F/`J&�귤=/RL��<���?���?����?A͟ЉU�M�>���`�/�eoL�i�dӚ�w��O����O@����$�ͦ��T��u�V��	6� }3u@�-([ݴԛ��-� �	ڰ 8h6-�� I�)��a�%O޺HN�ı�h�O���6�'�?��"���<���?��C�D�l�15�
b.h%31@��?����?�����Q�ݚuE����IڟL�f�
�c����C6'rH�,�l�^r�	��M��iۘO���7Cw�)@�,ҷ��0(���<)���2A3.x� ���L2"��Ȅ�yR�ӪH $��J(��q' W��?����?���?����o���D'�
a[�a��K��E�d=��'�Ot	lZlyn��I�(��4��'d��++C�hX�Bb
3f�d1D��*K�'DB�'_ā��i��i��?*d�d��M����%'Q >�*�
R Z�U�Z%�Ė'Db�'�"�'r�'����K�$�Zp[�� #Q-�`�$U�H"�4h�z���?�����<����]�� O�0jT(��	����m���S�;�mRQ`��Q~��!��^W�2�I1� L`�'2\�ÀEݟ01�|�V�H T�ӳ�X�$w�8UA�%�K8�{��v���z�O�����Ľa.��1�h�-$t���i�O��o�T�������I�<�_���C��s��Y4�W�Z֡oQ~dQ�_lb��Ӣ,��Oy󎈓`$�#3�֢5sx!�����Bhr�'&2�'��'"2�3Bd�"�'C�K�<mÒɉ1\����O �Đ���8f�KTyr�m�c�(*�e��jX u��'G7�1�A
b�	��M��iQ��#Μy�����XQ��K�Ǟl���']�ưi������'�LQ'��'�2�'!��'���'�U3Y�Uc�Y($�87�'�[�x�ٴ�v�K���?�����O[0���)��9htp��mE�,F���*O:��'9��'�ɧ���'�"}���52#4��"��(c)�}�b"R A��9 H�&:�	�?QQ�'$��%�TyC�!wo:-�d]nc��)�A�Ο\����p��̟8$?-�'6�7� �H2ĨK.80�#��C�6,�yP�*B��I��M#�2�>�%�i�2(�g L'.�����@g<�ic�
�m�8q�)og~"`L�,�Ӎ@-�Ӌz4�L�����C/`����-E�@�d�<�	�����J�}vx����[H��޴c@~}�-O��6��M������^q`�Q�h�i6�z�.��`��nӐ)&��&?�XFd_�m��y=j(p �`QV�s"È�y  |��'�b�f�'7��$���',2�'�Q�Pi�Jux��%O�����'��'�RQ��ݴj�4�b��?���PY�Y9�a �\<n�`��o��d��k�<����M{Ɠ|����=R]��-F�L"x09� ��?���vܺ����H�Ԉ/O���W �?�RCw�P��	��!y��e��>GP��Q��OF���O���O��}j�'�ntX��Ҡ)���w�L����[���P?v��I��M��r�O���ҧ\h�dC0D���L��S�'�7ڦ۴VC�P�ڴ���?<P�'9@���Ǔ'vP��v̐�b����-*��<���?����?���?QD��P`¤cײ���ke!>��'��7�H@�$�d�O:�d3�9O��Bw��3z�U�R	Ň%J��b�Fh}r�jӐul�4��Ş�*#'Z�V�� ʒ9d8p6�"r�q�*ONX��`���?��"��<�@��t�I�b�I�xO)7l��?���?����?a���٦����<)�E�1@�b��p$�?)�v�
�.ɟ��ܴ��'� �?S��h�N����.� ��q�Z 6ߒ����R�b���)i�t�Ɵ�
qa��Y��<�'�y��5uR����P0{�:��DG+�?����?��?���?i���˧E�	�D�>��3�J�d%�'A��h�f\���O��d�ަ!�<饃�#���"��D�0�6����	��"z���
1e��7�"?�KD7j���2�T�.g޹�vE��VC.����O|u�H>(O:���O<���O�`��H�.[
,�ya�T]�Z��%�O���<�5�i��lC��'���'���\�^\ې��7=����@�?E4�U��	)�M��i'�O����j�mR�:��	�0L܂o��۰���Rи,�/���D���L�O<xO>���+,��b�Ď�M~�`"ų�?Y���?)���?�M~�.OVMm��D40щR�`7l�� �)h.��1�ß���(�M���L�>	�i��g�H<R3�Z�X
f9zC�E�N���'|�&8q&�}�&�<�&8�sh��T9zɟа�&���P4jǢr_M�'i��H�	ӟ�������I[�4ײ<��:0EHH�~5ʧ̀?��QB�'�"��T�'��7�l��X�LH�u{��u�QPa��Ϧ	�ߴ(��']�OĠ�b�i[�d͓e��� ��<	��e�Tbуk�"�	�x2��	 Ld�'~�Iٟ��I�-�LQ5�ŀ4$Ș�,E�>�
M�	����I�L�'7� Qnl�D�O0�� =Н!+$LR��íQ�j�㟌˯O�mZ�M�x���!"| l�Q����x��K�[��0O'F��R&�9tVY&?͹��'{V]ϓWF�Yc"ᗭ� =薦��<�]�I����	ϟ��}�O��(LiJDHADM��x��$����aӠz��O������?��'8��(�#��(%�@�V�2��yq��d���o�3j�o�E~rnY#4�����WnF�M�$ZV��1��TAї|2\���	���䟼�I˟D[����V9�YY�eϪ-�
�&)?y"�i�`m'X�d��U�'C�	x�Eϸh�]Z��7.��-�4U�Đݴ%J�F�6��I;B~�eе 'g"J �`0�$IS�P�Z�˓SX~���$�OtY�L>�*O 5���.ö�f.Eb(P����O����O��d�O>���<�i��@���'�n P�iW�j�{�E��`7���'�V7�8�I����Sڦ��44�A
c;b P���zɑF)�<#9ݴ���%'�NiP�'���z�.w��Kqf٨t��rW�P_P���O����O�$�O��D3�'(��=�C��H2�, !ᎌ,m�u�	ßL�Ʌ�MS�E˲��$�I�<I�ߔI��"�a�)1�L�c6J���c�&�y�v�霭*��7�#?���
�&;�	��av<�2���9c���c�O�x@L>�,O�d�O���O\s���t��a91o·3�@!"�O��Ŀ<���i�����'���'n�ӟiN~&� �{6�k㈃g���4���)�M�ѷi<O�I��D\�eL֧lg )����4=��@مo����a|��˓�����O$L�M>��l\UY���D�I.��dD^��?���?A��?9M~�-O|�o�M��0ό%5~��h��& ��q�@�`yҥs�0��h�O��D@'?�|9z$%ݸ ^J@S�畚*i����O���1#h���Ӻ�&�_8���<R�nT>i3��5H�.mN 	�A�џ�'�b�'��'���'��5	v� �#��W�f�p��ۤ(zF�oںD<�a���L�IO�S���4�y�R(H��[P�D���f�\��?�������z<X��4�~" �* �����h̲4����ڊ�?�w���dZ������O�$5v?����2���#K(L�8�$�OX���O$�lɛ�LC]Q�I�k��{�k֡K�Pu����a�5��	���v�	<c4�J�� *�0�)L�	��L�'��q�l;
�&X�����-��p�"1O�8��+G ���l� ��Mr%�'��'�2�'6�>��S�? N���m�Zo�u�AF�����Q��'�$7�ɶ4���O��n�q��:�K���L��"��'�vu8�?���?i�~ݐ�ش������U���xY��ڕ�$X+�#۪'��d� �8�����Ol���O���O��D	�3�^�"�
b &Y��R�p`��/���a�R�'�b��d�'�����Ϋ6����%���@���>Q���?QL>�|:�B�=�����
9�%CKY@t��C�;��d�!qm9�`���O�?�<t�w�`��oԶv�u�q�R�?����?���?������צ�0 �̟[�j��IkL��iS�&G�%��̟��4��'�&��?)���y��R"Q�-��3pԉ��3D��L[�4��DHs�&)���E��*&и�k�)�pdr�JS&B���D�O��$�O����O��D.§rv�,�"[�iޱP�]<�\�	ӟ`����M�t�������¦��<Q@��&��� %\�9�>Ml �+�'5�6m�Q�S��HHo~E��>�8��צX�
�� �,|������L?iM>�(OX���O����O��DiZ7S��q�
�6O
`Q���O*�$�<��i�h�dY�d��@�d&�y������L�#�x �g�@0��F}rGl�(�m�>��S���=+ujp)v�O�s�t1Q5�-�޽�B2L��ӇX������M_r�>n���Q 0�jN�P\����MV�n��;�?Y�v��"��E^@q(O��nW��]�����Ms7��8V]�|h�#-I*Xr��_����k��Y��/v��T_bx����� X"ɟ�,���ܪ6��AcΗ2`\��F�'�����|�I��|����I^��,ҫl�g��j6��`#
��n�V/E�H�b�'gr���'d7�x�xb�刹`�ޭhd%*����uǅ榝ߴs(�'N�O?n���ij����,4�3i?7_p	pe�D�EM�ʂ<8����IW��'����$��"{���ը$y�l@c�J"a�zx�	ޟ��ן��'a�6-B�Q����O*�D�e"���m^������D"�.�"�dIf}�~�&�lڑ��R���R6q�����p|11��?��C�+���('V��dHj�_Q�	�v�:��M؛j�^��A�TF���O�D�O��D$�'�y�d�' �}a����%��� 1�B%aӨ�
�<���iW�O6��> c6��AHC	W��P�gÄl��dߦi3�4'�Cٱam�旟$P%O����d�w���buB1#)����
���'���'�r�'�2�'+B�'��l�D��-��Ta�#S�o�:R\����4-u�U���?y�����<Q	��
���r�O�g�tɓV�Z��	ٟ�o�6��S�S�K%��yaL�14��\ �h0+l.9ӦfU����'ǬL�d͛؟�g�|]�;Q�^,@��L�B���R�Ō�d�Iʟ,�	�P��ly"�u������Ol��̜�b��qط�	�)��t�Ы�O�o�x��v����M[��i���$�/J�:����6Kģ0��$䠄 ־i��	����g�O�:!%?�λJ��!�f���F���L2�
	�	ٟ���џ��I۟��IF�O��-�N�E!��Ey�Ȉ���?��>ț���848��'�b6m/�7���3���*�q�_X̸sԒx��f��mm��?��ENæ��'�\D�PeP�HW �a��o��/Eku�I6~�'m��ߟ��I��ə@{�8���}�~	'k�6_$��	ޟ��'�.7��~�����O��;�FC��]ND����iŘ-k׎Y|y�o�>Y�iQ�7Mn�)�d)ؙ8������;'�a�6��|�1r�/Q^�s(O"��ˌ�?5�)�.$�H���3j��L�%B�)P N���O����Ot�$!��<�P�i����ĥB4�}�$Ì�"���[�Q�]H�	�M���ì<I�t���'��'�X�`��۰]}�lK�4xA�� ٸ1F�&���".&����[b�4J�H�H�0B˧Z��@�ڢ�?�(O0���O*���OV�$�OR�Tmr� Ć�y0�k�ϮSҴ�4&��h,On�7���O��l�<�� ���D���K�e�"�Bc���M�i�O��,��W�aӌ�	 ~ MjwnR�+v�(�oE���M�4���D���?����d�Ol�䗣q LY���[��C���R���d�O��$�O��%z�F�H�Y�b�'��EJ�00��1�L_3D�bJ�J�0�|��'�j��?��4d3�'椁�%6M<>���L��+��	)+O<�(�gI�1��%��%�	�-�?!��l�T��C'
��)B7�ɚJIx��O����O>���Od�}*�'}>��pȋy?�ԢfHY�(��A�� ���ʇ�_�"�':�6m�O\�O��i�z�4|zD��%	#|a�VfL;��D�OF���O���� d�D�E*T揂���K^�r��٢c��1�*����ǻ8�`�O.˓�?���?)��?�eV&��rGW�}U�-#t�!����,O��m�S|�I�t��|���8|�c(����}[�AL��@D�4\���ݴU�6�8��	
�yd{�K��=�T�)�O�FA2�y�N6K��˓fx*)0f�O�ZL>9(O�sg�+z�
g�?���YBB�O����ON�$�O��Ĺ<�U�i��<0��'�6�j6�� ���i��5׀�ڡ�'a^6�5�Ƀ���Ц��4y�Ÿj�8� 6�K�LKr��C/i&8�bݴ���W!��a#��B: ���睎: G� s�N$Z�,�.�����O��d�O����O��D!�g�? ��P�լX�j���%�_*��V�'��'H`6�M%߬�'D%�6�
�����w�Ļ1��Uo�<��OznZ�M��' �	��4��DWP�[�M��WGj!+�� (D�r'Oָ�?�u�>��<����?A���?� �N�Ez��c/c}JyJQʬ�?������5�����H����O�Ry2'���d��V �И#,O���'`~7�\馹�N<���Д��K6�\i&�@�!�p����M������h���?i���'W�M%�|����6'p�L�Cmԑuy�����{����ٴu$��7 �DE�X>����<&$�����?9�i��O��',��.��js ��7��eh�cۑ(B�'F� �3�i��?�k3aP�?MhEW�̢�/�)w��W�0#;ĭ���T̟H�'�a|�%[9�p="$�ָqz /F�ms�F�ңB������
#�i��䆸E���t�(O�fł���31l6-��bH<��'���)�H9 �4�y������	ԣ6�HQ�E &���K�@ <|�I�XO�'#�S~R���5&�l)j��@�� ��I��O�<lZ�P0�I蟄��m�-&��zX�	��?k9^U�?�d\�� ޴}��F0�d���A��%���14ǁ�r��˓��՚�k��M������k?�'X\@#q���l���Cg-����Y�'ozy��#�9,�E�F`���� ��� ����m���'y�6�)���?5�ҦĔˮ���
�tX؋(�ן��	��	�!��oN~Zw.X��v�OgJ��T�/!pȼ�ædET��dd�}�INyb�'���'��'���Z/,P�2���(����N3 ��Ʉ�Mc����?a���?AH~�!�� q�^��Q�e��n�� ]�px�4
כ�:���ީED@	H�
�a�8�Z��T�J����� f��ʓ@v��U��O�݊H>�-O �Q$�H(T ��Zyn}��B�O��D�O��d�O2���<��i���q�9Oi����S蝲a� �D�FdC��'O 7�#�I���O@6���y�*���M
b��k����B��7�2?Y��v��Ǣ��'�ygI�G���V)j�9����?q���?���?����?9��鉩�❑E�T�^���rc�Ҝ?���'M��{�4QZ��<Qq�i�1OV�XRE�"��蒇�H>Cڶ@I�"%�SѦ�ڴ��"���M{�'z�b�%K��{�A�rdv��&Ή[vM1(��|!��|"X����П��I�(��a��F�Tɻ�$�*o�`I���d�Iyy�t�(`c�O��d�O��'tN6q���&s4@T��F�i�'b��)���M}Ӿ@&��OyH��T"]�	:�t+�.	�j�J��?q�VY"� �'�����Aj���.�O�!��a�1�`�؅ �'(�ڱ	�O��$�Ov���OB���\�v"��c{���Ƞ2����G��:?��+�W��S�4��'����������l��B<[U8Q�ǁ3}�N6MXߦ5*��]��͓�?���^���)Z���d[�QY�����Θ`ԮM![��$�<i��?���?)��?�ʟ�ACf�7c�V�;��{��MZS'x�ڨ0G��O*���O֒�����͓W5�d(��εs���CN]"xLpݴ,�F�<��(����P�6m��|js�[q3.D*ZG�6	�a��únZ�
�d �4�'���%�$�'|��'�yHG'���m��cғ���&�'kb�''�Y���4_�FL*���?Y��4�f 9t)S�74���@Ǐ�r�����>9g�ij6-�]�ɡ5�b-؃���zSd#��|�D��'T��P �:p��u�U���/Y��`��>O�����A|�Wσx(��'J��'���'n�>�rGJ!��I�)E�ܩK�`��5c��I�M{�H9��d��E��s�I�?EXdH�"��X��MR�}k��C7��蟨�ش���,��x#үd�^�ݟL��_�u��4H8ki�4�pc�-C�ؐ��Y:U�&�&�Ȕ'�"�'���'�b�'!�F�
��� G�_�n@��Z��k�4G9�����?A����<Q��ۨ�XĆU������#}���O��m�����O�)�<>��-Zq,�l�|�6��)F1hG����@�'^�e��ܟ㳑|"Q�hP�"�4*��\�FkY5)6	��M̟����h�I۟��	gy2ho�
�BC��O:���qy*,q�!жS��`;�N�O�)mZF��UZ�I8�M���iX���qPz1��˟�)ɠ%�7doT����i�ɑm޼���O�,�'?�λxJ,�1鋱�B������,�I�����z�O��
�	��n�s�&�E 4����?���JB�&#@76���M��yr�I�Go�ب"�Ĉk��d��(M<òi��7-䟪Y0v�{�������$�ǢH�����0�v���fK8Z�r��X����d�O����OT���8D�zA�+�$0�vݲE�508\�$�O�ʓ1���B3T���'�2�?�"B,��nAV��.�����Ǫ�<)bZ���ݴ"���?�4�����3yd(fÞ:5Xi@IKy����g\A�(i���<��'W\h�����V��A� �(�$��I\��5����?I��?���'��$��� �*�l���u$C�"+����R0���	���ڴ���?�PT�t۴]$�@"�%�|i ��.^��4�Q�iK�7Ĳ[A@7�4?q2N���t�}��ό7l�ջ��ӄLԆ]�f��?�.O0���O����O����O�g�? ��x�'^0A�pp�2H�W���z�Dn�>��h�O���O����$��A͓8P��rb M�9���z$�B�a�y��4mO��-.��'�i�%06͸����4SD¥mQ>=0h`�!
�OfASƠ� �?��/���<����?9ׯ���d�`.,�Š�#��?a���?i�����-9��۟��	ȟ�����	+����Q�5��"c�I��wt�	��M�5�i^�O؍�0��:̜�RR-�R��,0I�<I2�5�Z�2�`#���V����y��	SR��цҤ�f���?���?!��?�����,��kψ}�<m�"K#*[8D�%�'��6탧q"RʓBV�6�d��F�X@�+1Xy�a��e!� a6��O`�n��Mc�i���Z6�i��ɂ�@	��O��u�hh�B��T���(�O��ey��'��'�B�'�fW%,�4�٥��To�|�łM�C�ɀ�M[��/�?!���?�H~�CH�	[pO:V$r���#��}��Z�U��(ٴk?��4�4���I����il�v�(��"P�td{�C[2`�v1B�Ȼ<�m��bȌ��������R�H�ɥ��A�N�(�/�~~&���O����O���O,˓F���U1>�r	 ��4�� ��^���9�j�2���o���q�O�m�M�$�'��@
�{f<���9B!�A���MK�'��)�[�B�SJg�I�?�;D��$N�&u��JƨB�v�j��	��<���<��ӟ(��o�O�U��b�e�1��ƖX�H�����?9��ED�(�P��'�d7m0�Dw+1������;�`=0%�<W\�O��d�O
��m�6y���'m1�����\N��Y�hʤU��j��
�?���5���<i��?����?i�a�D���3Q�q�B�#麜�I��0�'g�6�1����O,��.�%��Q*�W%L�#� �r�����������צ�ݴw#���ӮG�n����H%�4|�4	\�+g��Pi�E���y�<��Oa�DI����|�b�o] :��&�@�21 ���?���?����䧂�����Y�M�M�p�.�x6�p��
%�,��ޟ�ش��'��uI���S
\��#��
I�Y���^"�:7����i����1�'�p��d��?=��?-b��L�6^y)��F/Gn�0q��O���?q���?���?i���I[�w�Za���{w-�Ac`��7�W+�����Op��:����M��'^�I��=>�����N?Ǽ@�ѵi	�6��r�I�?a�S�?-�T���5Γ$' ���`¬�Z����K���hr��*�Rp,�O�t�M>y(O~���O��á(Ån�v��s �}6�Z���O��$�O��$�<��i�`�h��'���'If�S�@D(|*Ha` � !��UYC�|��'����?�������5Sag� 8N��� ��\��)O��gΜ"�*�"�K/�i��?q�kf��㊐ 8J����]]�DC���O����O����O��}��'���觯1	��q.S�.��\���rӛf
ح{!�&�M#�B�O�$��v���
����'�K!P�4 0O��~�bqm�o}4Xn�q~b�K�!N�,��mV(Cr��&`�}�Y�d�E������$�O����O8���O��D�.���Ru��dnx�g�ܮ|��'���[2b�b�'\r�O6�s��(��Bu��1c�ɗgN��q��������9b�45�����O/�4M'� �ME�&1��Q�(N?^����<��I�:�p��'%�h'���'ۨhy���
�8�DK4:�iX��'IB�'z�'�2P���۴P�D�����)��X� ��bC�a徵�;�F���J}/dӆ�oZ��?1ՎE�i�ʼ{g
�<�4i�GK��O��m^~ҡ�aN��Ӡ2��O~�ND=F)�1Ř�5~F]��X�w��'s��'>2�'r�ӭv����[�d]�f+��]G����O��dSԦE7��Wy�o�0c�t�1^,p������L�c��G�	��M3��iL��,)����,� E�;2��SLJ�5�VG�3���(P�'�:%���'G��'s��'��� ^=���e�ג�8��G�'��R����4͢����?y���	�W�&�bc��Z{ԛA�`�剗���ަi	�4^�����M˶��s����N_69r����W �.���<i�'P4���"��PW�[��5a��X���7����?A��?���䧷�$�ߦ�B�N��%���N�4�f �(䈕'"x6�1�	����ʦ	��/ �P�U�E){�X[bF��M�%�i�j���iH��.�R�5�Oz�p�O�I�0'C�<���ḃu��ͱ����O~�d�O����O���>��GΉz���h�:@�\�f*��M[A����?i��?I~r��\Ǜf2O�D05A'T�!8P�	<~Ӣ���nӦ�lZ�ē��E�>Ds�4�~2"�W�2�� d�Xhؽ�&�8�?Q5i�-C���e��@yr�'�B��G�.u:Bc�p�a���K"���'z��'��	)�M�0�Ǻ�?��?���J���*��\#`�R*0j����'kf��?)���J(8��䡘#\��Q��7ag�A(Ot�[D���O�1�@)��	�?a�``��S��Ƣq�d�
��Iq�O��d�O^���O|�}��'08��$F/c�������
U^�"��a��l̮2Sb�'g@6�!�I�?1`�k�O�@I�姜Sv6h���H��ܟ��	�F|�Ll�U~Zw,6Ux��O��h��\�#mF�I]i�n�w�Y�w�>u�Ѧ�M��Sx�6�bL~�=� ̨д�I�1��XCc SB�]��"O�y�'H�m�$@ &��`9P����ل&v�pI� Xt*��V�G4������~�t�`�$��t  r�ފ:N�akĮ�T�x%�����jhe(K��aJŢ�=T��[s�r�`CK�j�:a�7�R>Ѐx�%�lQ�6���~��ya\'i�$
����u��	�I����r�/J�z��h�e�j��X8�	Y-}����&㌋M��[!�APR��Y�����$���iWf����ey��L�f�P��ر��g�q�mH9˒\�A�i���f�0Ǿ�0�˞	=܈��^�s*��S1oM%��9�B�A�!��ɚ%pOR�Z�M�$���b�l9n�t	���ש|�$�2h p�N@CW̑/dgM��H�8��Q�Go3z�$�[a$�{�l�C&N��x��Ȇ%+8���C���e��ҟ��I�?��O��].��gB�A5���ޙ���3��`�$�!�����O��k�N�^ ���;��:FC������ʟ$�	&aH|(��O\ʓ�?I�'��#�j��&b�$����l�� P43��'2�'�R"�	�
q�	ڥma�F �0~���'k"a����>�.O��D1��.=�z��pN\=XP�8��ю�L�������O��$�OJʓdDy E�,P�.88��X���ꆥE�cS��xy��'��'���'W�,���>q9�Y�
�\ �dɱk�'���'Q�P��zsR�|���P!"ܲ�l�=K숫#�ǟ�������p�����2 q̓GS:,0fcXCRԚg��� ��'!��'�"P��9�M@����O"�ϖF�yhbc	�
$������O��=���O��d�",qO\@ic��;&���L�s(��!��'o"�'����&���]?i�Iʟ���>�T<*�Ո.��q7�� �>�'�t���*E�!���t�ҷ1lj��0`��D��ų����?+O��K�������ٟ@�I�?�ٮO�B�O�I�g��^���*�`�O���Oܪ�N�OD�O~b>U� �ELa ���L��c'�Ot�Y���Ʀe�	������?=èO�˓'���1���dx����c�����+�F\A�"���Od���II
]�L4�4��B�O��$�O���;&���?Y���?��'�l9ct�ׇ7G������B[�FxBG��g��'+�'��A	"2�d؆���E�\l��]�L�2�'��	���>.O���-�DF�:��\id����K��˔s4x˓trД�J>���?����򤂹C_�:��S�b�����HI��BP�<I��?���䓠?������)J�p�/B($҂�� �V����?	��?�,OxLr�b>y�Ul6I!roD�GZ�Q��OR���OD��1���OF��Z-(����B������9,-|�s��)v��?���?Y,OF��v�
�ӰJX�H��T�M��� N-c�"$��ڟh'� �'�H���'��(1H%��Z	�,t� �ҖBu����O���<aC��1J�O�3��\rF�B�h�z�T�,V��U�V�|B^�X��ҟ�'?�	��� ���#~m؍����_�tE��Myҳf~<�ݴ���OB��oyҧZ& �9�T�4j�u�䙻�?	(O����O����� dY��7;���é�i!�����O$�r�^秊�I������?y�M<�'g�
���Qxp�a`��f�#�K��E{���?a.Oh����<P$�U�Z�1���p�����'Or�'b�蘑9}�)Z�O�l�!c��l\=�T�^�v!x�p�h�'�d��t�'T��'3\����	!LиYXA� >	���'¤���O��O>�O$:��aD$A�J)rN���-�<j�4�?QH>�����O��d
���f��R�ϳ?�0����
����?�����'���'�J�+�
����NS�PĘ��=�~�[�y��'��	��Ļa*��|b�(�/tC� �1"�'o�h1��������ӟ|�?y��?qq͕2��*E)�Vf<kA���hL� �N�����O����O�˓xu
!�A���
��B�֝�VND	C�R���$�4L���'��'��ɞp�\��	X���*p�XA�'��\�0D�i��?1���$�O���*�|��?��w�^�)3��&f��#��I�A�|��M>)��?�J�
M�B%�<�'\�����<�^�����+��@��xyb��>wb:6�|���R�Q��!��/S�\8�4��CX舑 h�O�ʓT�.�������'#/�!3сL4����$V�=����m����?	��?1�'��?���!�TY��	]������
ٟ���S� b.b�"|2��N�\P�b��M�"�k�"VB�ԍ��i��'��!��t�FO�	�O`��7`�N� ��Y=ZÆ��#F�`�n�D�O��$"��,���ǟ4ϓy���y�oQ��
��ݗP�b�	ܟd�Х ky�]>a�?�SE�,.a�]�$*�+��8y2���To��'^��'��T� ���,Qb����LG֑I��٢1lm	M<1���?�*Oz��<���vt^�`S"�`AnQ���&�?�����?�,O��$�;���Ӄ9��aR�\����i�/	<V���O���6������I��NP����b���`�b�=c���
P/k�L�'���'�"P�"P�і��I�OLpӇ�R8GC��1��F<?f�[��O���<����?���#�����$��6�2<��n��sT�X�5Q2�'�RP�p�������O���4� 4���G�h�u��Y�����W��	����Ɋh�	⟈�I���'T��w@J�8q)��� m�4�	`y�5q�7m�O���O
�)�v}�� �A�!h�a�����t���'����?�y�\����X�'4�: ���*���x��QA� @�I#\U�`9�4�?����?��'P�I]y�_�Z��I�wJ�@f�0B��W�ie��=�y��'Y��'���$�e�d� e�-Ўt��ß�j��m�ϟ ��џhQ3
���d�<����y�.�!����
R
�c��%�?�����#z�\�����Of�d2:����
N����R?x2���O���`}}"Y�T�	@y29���I+�X8hgO�R�J(��X�41t�4�I⟐�Iß��	cy�N�>��QCE�	�h���� ���>�-OL��<����?9��S����aK�3��C"�P���ID&N�<���?a��?����$�Af���x�*��B��/m��ag*A���O:ʓ�?�(O8���OT�d����DC���߈UP��mM&	�˓�?y���?�.O�����u��'���P��-浚�m
�j,}S��'tQ���ڟ�������	A~���T��#��3g���=�?Q���?)O&l�� HF���'#r�O����r��6�A�&�7��a1vW����ڟ��������n>���>�F5 ��L�x���O�ʓOhm��i\��'���On�2�
e�gi		V��i)��>�f����?i�\b����9O�b>��U�Q3$�HL��Z!^�H��B�O�=�+���ҟ��I�?E��O��Zg�1foL8I(���ƿdNTQ������'��Iq�'�?��ۧH�=*e�Nb�P�H���9ɛ&�'�R�'�&� �H�>)-Ox�s�Ј�#�F�$a3�kL�f��fk$���4Ӣc�d�	���	�z8&P8$�C� �@��9/��IşP3� >��$�<�����a�if��?>n���F&�*!��M�<����<����?���?	���S�|�X񧏗9Y� �Ꭷpv4�d�T@}RP���ImyB�'v��'� U v��;a��b�o�QkzErVO���y"V�H�I�����Xy��b��IN�l��X2� ׫�XQ��n]���^�\��y��'b�'b!�'�R!��l�0�Д��L�
����S�p�Iٟ �	Oy"�[��꧛?I���/`�i���Ab�A��%�?�����$�O����O��z�0O�˧{�[�U�6�dE+#ҁo�H�Z���?I����H. ���Ol��'R�����%E��,^�'G���c39"�	��	ϟ���Mh���y2�䨳
Т98�P��%$1�e��'��	���4�?A��?A�'��	(K0�Ǧ?K3Z 0�Ǘ 	��������I>���Iџ�'1�2yb/��O`� sħU!w|���'�d�mӾ���O�����ܼ�'w�I3�H�2�]<
a�������IU(�Iן�'��4���5��P�F�Y?����V<���l�؟(��ҟ���ۃ��D�<)��yZ(��6	�9]��`�!ǫa������?�-OBH,"���O~��f>5�s�SQؚ� d_�D���R��O8�$+EJh�']�	Ο@�'\���}�ѡ�o� ���4C�I���~y�'	B�'��	a�"Fo�a�$�Hq퓺 ̴`���ē�?a�����?i�~��)��62�=B��� ��Ԓ����?q+O���O>��<i���/m�d$L�0e8��O�
Xz��m4���?1L>���?)�
��?)cc�N_�y�3!�57����#H����D�O����OLʓ}�t3t���	ޜ�|a���%��l��ǟ8H��';�'��'	�ɑ�'z�Ic5�`���)>��TyD	��;oP���O����<	1LɏDۉO���Oq�8�*� х��8>L�(�7�|��'M2��	�yґ|�O�R���&� ����"��X������d�o�J�4�'��D�<�0o�����j�Z�C���G�Ο��Iퟰ8"�i��$�P�|R�K�0X���'b_ `�� ����,1F�X:�M����?����p�xb�'����o�6�����)�'A�kr�'���'��'�����"�$"�.�� �j|C�,|�t%n�ǟ��I̟0y������?i���y"�� �>A�ǃ_ΉR�����'�Q��|��'&��'�u��@K�#��}��l!��c�'B�"(7b�T��Iyr2�@����L)��]�MY�9�V��8�at�`�'�"�'%�O���ҋ�6Z�&Ɲ0 �	�7A�)Enc���	U��������/#���lIS�2����I�&�)�����h�'2��'��Q�V��L���iƇx�\eePJ�;V�O�Iԟ��IL�	ԟ��	�hX�4��5>ȾQh!.�]\>$�bϘ�OcZ��'T��'.�^�����B��'	���hA�W#4�,yQ��F�7 ��z��?�K>q���?�7ז�?i�O`�01�_��悙5�t�H(S0�?����?Q+O��R�b���̻-�t�VK]0d5��@T��?���)Vi����Sb N[�l�� H�0i:��7��ȟ��'JĐ��A���'�?���y��7"�l�����e˘�4l����ʓ�?1��0�?�������..����b�3TT�����!Tc��ح)��6m�OV�D�O���[}Z��� �l� `_p�`�0d��x��-���'S^Q�'G�X��2��&pu�5���h�6�
�O�����4�i���'���I sh������O��nm����Ԕ,���@�ɖ`����OL���O�(�P�+�i�Ov�D�O�m�W��~��yU-�y�ưQ#�O����/��\�'��	ɟ�'����w�!W��I^���o�b���!<���y��'��'��� 
~0m��/��*�jș��X�PN�$�vOҘ��D�<A���d�O��$�O���ǈ�QFE�2S܁�F��N�1O��$�O���<Q,�?2��D-F�\��i��1�l,򕀙��?1(O���<9��?��O�Ru̓ I��ƮDD���O. ���?���?�����	-	L�ON�E��E�W� �W{0z���S�'����d�I�좄�w��O�t���3�"�I dU�
�>���'ub�'C�I5Mfn@�������O��	�J+����HV�%�K'�.˓�?���?Qr�T�<O>��O
�801.���j��d�ɡ2H��*O8�D�o�|���OZ��O����O��Ӿp(̜�@`�?�y�g��(�����O��$�!)E�uq�����S4�<9g�ۓ�t�v/R#c�RǲvG�7�O����O���Ww���� `$#B�#�l���ē�l�����L��ԩ$:���O�2��(V�����HF�x@�Ӫ?�h6��OX���O0m{QG�M�Iğ��I�<	Տ�$r֬��1^=C�j��ӂ�S��p�De�?�n(I_R���P;8(�IC1gʌ� ��5p(��0�@�}�<0Fm
+����&�? *b�'�2�'fM��j�^���%]�1a��Ke
��l�
�Qq Z�y��'�r�'&��|�<��P��U�@���'b�	X��L#��i�b�O���O�D)�d�O\�H�jM���+3nA�U�fh1�ߚ<:0�W#���^�h��1)@�p<qS(LH�,0�������R���F؟����Py|�͒�!�5a�
�\̢m{U��2z�Y{NU���*�ݻMQD��FΕ�=�|�P���H������$VG�LQ�f�ɰ�h�c^%�e�O��h wL�!����'fV{o��z�li�2j�wv�� �gæa�(�
;�j��0���Bb� ��-�O���O���U�?� �d�OP�*u�Ɋ@��2}�U�шr1S"a�f���΅1�vUi��=?H��D~2nɨ@APA�֭�klv`�´d;�l�ā�Զm�%@���6�
���m���'~�����M�Ώ�a�w�ڀ|lD�� �ўxG~�̚���<(r��k(��:7���%Ȣ�,���µ�l��A��	ty���)7��?���\���P�C�i��(A��P5ri�(����4�I��~(k󎕺-c���.�8�?�O~Α��\i&|;dI]�`�������/&rb����+�M��	ɞp�Ո��L�I6n���HO��V�'}b�I�/��xv@Yp�z��7L�,��d'�O�X�狏��D�S�g����'�`�'C�y`�֐�4�I�P����'�"��w��>�����	�3�t�$�Or7́!����@7*M�p)��#�X3��+Zph�8w���;���S���iG�顆#��@���&V쒽�4�� �i�E��t���)$"�?7�L�/��x#� �,�69� �F%��E�?q�����ԘxB�� z�����O2J��-2$&�y�ZN�����ShdX�CD܃�(O:�Gz*����e��;a���"D�o�ٻ�G�ȟ���!i����EE�������\����uw�'q�& ��W�4�
J_,d�>a��L�	k����?�&y3�/>5
p�������(�6b�l�r�l˰+��TJ@�+�B.˳#�j�Á*J76��g�'��rs%��}���A3���x�Or�[G�'�"�IT}��F���������yH2���y�Q dh�r�Vv���ᤞ� ���EzʟZ�'���S@�18�L��ΐ�g�YKF`�v�84���?����?� ��1�?�����4��>������13ڡ	$�Vӆ���R���"`@J� ����՚d��e#��F�dd\�6'�4u�ibǋ��k(���gWpu�	ϓ^����Ǧ�Y&��K*�z��C�?�����E)D��$��'-���h�*'�����N'D��*f�)4�ԘG�8:d*��񋯟\��}��g��6�O����~��%F�Н�7�D�v��0�P!�޵2�'Ir�'��yp���0S����H$B*�T?����g`��Sg�&d��G�*ғ92�	�� ��l��i��S�]֕�q�&�u�1�։s60"=��!C���D�$B#�z(����q9�����>�y�N0�^ERC�L3)^��d�E�p>���>�҉�P"�ICB�QS�1"�$�h?��Za���'V�\>�Pe����I���S��/3�	)�+�:tz�c�8����1���k��ЧO�h�禝�u��\1j�ӗ��4d�� pӀE��-F%R��\!K�"~nڣN��4���{N �h_;m��6�F2���s�>�!�C^g�L�V �g��A0"O� � (�%9wP!�4�I Z��%!剽�HO�H�F�� �^X �cs!��_�Y��?9��Q<O��`���?����?Qc��j��w��S�D�?��@����O�@��f�rWN��D߸%8F�����%8�̘%�] 
m��$3���9��q���z`�ӀQb�1B� ^�f6�)�I�>)��ӟ��ɎS����*�0]	��ceB&�B�I�h(���v$+�rh�3BT�$sq�)�'-eT����͒u����ߟ�dٗ&Դf��Q��?A���?ɱh͒�?A�����ٯ.�2,yĉ�b��葁Fl�T�	��p3@���y��Y�;�DpiPF��c\JІ��4�(��VI�FX�3
�yrB���?ܴ�P,3�s�U�ʛXԹ�d\i�<��.W��ؼ{��ACTT�cbIz�<�0�P%G��HXP,ַq_�-Y���_?���$Xb���l���	O���'��`5�S�1\�Ȉ��a�Xl#Т�O*���ONhi���h<.j��S��
�6Ɋ��#Ҋ�R�A��HO�c�i��Q�SK�;%�V`����I=R6U��!8 �%���ɬm��$:�'!"\�t(M98)�@����p����)�Y(U:ch��BVa��F�f8��J�<آc1j=�� ���*h��뱟���U�M���?a(����(�O��dg��ap2�!c0e���*2��l�F��lƁ�	V�S���G��-&��k��v�LL
ר��MkEC�E�������Fgj�xA!�+r	$(�AD��M���L̟x�<E��4Q��px��V;z�@�6e�!5�D]�ȓ1�KM�D�����9��z'�"�����'p��41�!��E& �	��V�[n��'O�F�.{� ����'���'��f�����b�:q'��2����M3*�i��X��V�U�{¡	��rG�����Y5#E���$] T��h:�;���k�-�8N���A���09�'n�q����=��f��qì�s���*Ē1����j�<y�BJ�o��=��́�-u�$*�@��'�Z#=E��O�*,�� �I_LԐ2ն��T�����?����?��,��?����t)Y��?Qݴ&O���� 4��"ܦ'R�q���)z#l�?4pP q%�8Ѩ��#�ף�zQ����E���c�}��	V�iH���M��W$@��p"OT���T�.߈ �ˋ�� �e"OPa�&�3h�c�ͅ�C[�LrA�O�e�>y����l���'aR\?���)Z��-�2�Y��xX��[�����?��9r�A!�͕?g�@��'s���P�G�a�n9��f�3��"=)��x�F�:v��)c�PL�/Fh8l�G�њZ�T�˰LKB;&q:%IK!na��<��ʟD�I��M������ډED�EIʹO�8���'�6[���I�'����'�f���b��vPT�u �;/i^�K����m}�n6�̔RUV����̙y��&���zf�ݴҎ��#�i���'�2�O��5*��'.2�i��ai�ɒ�a.�HU�K���뒭�A���1�|�?��퓉?l�#�E1t[���ʅצaK2/�S��M�)+��08B��¬K��OΦy`�Ozb�"~nZ&!auPN�#r���7[�#�lB�I=~,t�f�	J	,�	��	EZ�<���|bg�֋q�.���̪QP���Βv~2�'����&���Z���'���'V�֝���.�_�z�G��!L`\�B�+^��	
��a#J��z��b�ʤsB�N9v��-�6U�Se�MA!4��T��	\���g�'-�U95΍'a�ۖ�k�t;�O(	��'�a{b�T�/����rN�XT�m�E�(�yRm��BR��j6�M'��ہh�6��Fz���M�S�*�+��Y�/�j`�d�طVA�ȚK���$�O����O\h	���OX�Dr>��5,���Dm�Ӈ��˒�Z@�_�G�PkAN�*)�d��.ð< >�Grȉ�v<r$ �g5r�@�U˕?�8P'`H�j )P`�w
T�P2�Ix"��yӠ�D,1q��)��&@5�X	
ɟ�?����'�2H��L� ��m��i��fu��'��` 6C�,30����*	};��x�'͚����"�1oџ@��M�J�=?Rd�7-]-~D�E8��'.��@+�%�O���OJa�,�M�s 0M��I���Ϧ�':���
�Ν�\!N9i�F�FYEzB.��M�2xE��ȅ`
R�tNۅ����	�$'�p��#ۃ�HO�:��'q�>�؁�4W�(F?<�^9�j5D�|�3)�#a>�`��Hאp̊��B�/�O<̤O� ^d�I�2���� U�B;tQ���OF�� 禩��ß8�O�t���'��i��1
����{�n�(��F	���9v�2'���&�|�?�e+@�� �*�;zZ�Q����q�$-�S��M����M�:�0���k��8�T��립����O�c�"~nZ�h��&@w���ӲVB�N�J�چR6�c�5M��<)C�|��5<$`H)���bx�9;�'0{"�'7����N�&y��'Dr�'~�֝ܟ���3F��!����10�M���?�0���@T���A�O �.�Դ�"�
���Kn�����/���S�g|�d�:׉�5��I�=����5lO�a�w���0��'�P�`�	��!��V�\�D�D-�:?����J��n�0����	��}�!늋Z��@����ȸƂށ;�����ҟ$����L�����$�O�Mjb)�&Yw�L��Λ/m��Ir�%\�M
��c���~A�5엾W+����� 2Q��å�/!����v��6If�g�Gp���旔zלdi��H�.HQ��*mQ��ڦ��O�7���CAlـ� <t����5BW�M���h�4�?�/O��d�O��$>�ӕ7L�$֨`��]��Nĳ%�C�	 ��Yq�Srz��+&M֢&~����M��i��'+"�''���y�jL3
� ��K�0U=�y��'����Ō�7B���G1d����:[æ@[K(]�n�C��G��!0OO���B9.]�I�l��yb%L"�f5*�	Z�*�,�C��	)�y�L�m�9ۂ.�:/�X@뜂�yүǶT�ֱp�΋>�p�)6ꓲ�y��  X�}�`��O?T�5%H��y2g� �q�U�\?��X�Ճ���y�l��7� ���,Y�a��Y��BW��yr�<n� �:g][����G�D��y���R� q�E�;]]gD��yj\�3���4�5]�	'�ɗ�y�+Ʉq[��@�e[ �2���A��y�D�z�z�f���&��&�U��y��ƨe�x ���G+��+�y�������%�;K�!���A��y�"l�*�ر���8�	F3�y�G�P+2���!�>॥��y2�P�a���BԬ7-��Kp퉐�y"F�2�<1A�j�;S���R�Y��y���*mj�lW4A�D)��
��y"D�s�uA���<�,��6k��y��1���P��7A�R�k	��yR�[$J,��J$�+V#�)5���y�\/!0i*3g]�L���aڮ�y�a͸@k�<�����A�n�yQރ�y�␝1�<3�/uY��E)����'�.5���Oid�Ҭ�]F�:AƸNюъ�'@XU�� ����G�)��	�r$� W�qO uE��O��A$�F����RCC!~Z��;!"O�C�I}���� �	%9�!e�i�8���px�Hju��3Br�dJ��Z�|�����%lO~EfO���$C�i4<u#��N��p���N�S�!�Q�#�^��S@�����Ħϼ.��O(����ʥ���dHA4(B����Rb�}�"O�����E�<��D�/3g"0�i��*�ӌ�Y����K�i�(e�0�'v�,i	-D�8�4�#S�8e�cfS8F�V���M�O�<%�3�O�G�G9�(�����E�M��%7D���F�).��Xs��As��#c2D���«!LD����<Q#�X��%$D����E���4*�a��� ��J$D�lbt�B��V�cL:Gf�L��&D�6K�KDl�a;b���i�Q�<QEg]��H����r���r�AJ�<���͸ <-P�.~�81����F�<� �ih�.8 � �*��� ւ�p�"Oh��Qb�͡��n��Ȩ6"O�D(�J	���P9�KHj�l���"OB���T1}�,@K 	�?�D���"O�,��
A6+)h�ە(-<!���7"O�L2��δ�y�6�΄`�(��e"O����Eb�X�c�	Y�`-�"Oмj�P�U��X"�"SX��A "Ol p�O�7V@�Vہ27p�!�|B-�26rb��>��s��(��Y���84-���0D��a5�\�;ֺ���ᅛXZ�yC�/�V�'��$㦮�X�g�W�B&��%�$�@�J�%)^�����~T�<r2
�:R���aJAq*�����"%���;U�O\x� �oՖw1������;B�q���*�x����qf�/]�`�	��SN���͢o&���0���ۅ��y%âܘy�L�Lf�qE�؄�~Ҍ 'e��PR�*q�.���A1�'k��Q{�
11�����;���	wx7i5B�N�qH�n>�!�G��q��6��0:��Ƴ��3�Ƀ&([�ρ�,g�MB���#WJ��� *�(yq�R�`�d*�ˮe븡(��5�:�@A��a���J��'� �ee6���{en2ШHh3(��XT���>���V�7v�#s�;T�X�b��|j3Ă>x�T�� csށ�3 ӬȰ<Y����j�K����a����K�S�8��O:	���X��35d�#��3�'NY���E �&N�0ѳ6Mٝ��L�K�d�7�Z38ՉT�O,�Dˌ?ET.�[�tM��r�K3B���Kte��V'�)$�#��i�U��V�)z�`ˌ(� �3�+�m�~)�b��W!9ӌ�@��ܴ9ф�pR�� C7lA�7���j�� [rĔ(;���#�{XLܒ��˲$Faz�kK<=�T�e�͐�v���B#V� 	�O[a�%� PC�_h�4ᨆ�?#v,Rul����K�m� Ւ`�� ~��H�4 �D~2��@���%��$��)������xs�n�.V2�r�ZB��pj�E�O���1�ð)M�uI�hʥCW�`S�.�n�OCj,a�91*�x�ì_���xɷ�>�GY�.PE��?��ٿ( HmѲO�Ԙp�9}6"�����Y�n��������WC 5ە��n��݈P�A����y� l<D�aV�V=�tg�����A1�N�I]���#b*�1O���s��.�R�
�O��@�nIĉ�ab��d�T�|l֐E���M�a��3\Je�K|���@6>)�l��DuPy�Ν�io�9CC'n�T��F��L
��"����O&�}�Ǆ���P���.��$Fl��'M,D�����:�b1cB�>��a��]|Г�6�"
Y�=�����L�7~[.p���OH����M�gE���A�=l|���l�7��%|�:�2J�H�� ��*Ml�h��M�`�'�>�"1���:���0y�e"�\t��?+�9 & Ym��:U�������?�֮�Q�v��q�9'�%�>qwCܷ"tNl#���P��B� K�U���H1$p4$�"Ɣ��ФϮ
��P�s��@��|��Kz��� .�'8���L���%��Lv]cuhRZ���~�;�#Z	9mV9�£�
"x��Fb̐�i&�Aը��+��*"�00P�bC>a�	��,�5[p�牃-&p��f���v\�OXD� ��1��O�t�գ�c���5��/86V,}��T�xnz�頁?��O����S!�=�|���%��1���N�gsPd*����gqXp��E��0<aS�("�t� v�)tl|(�!�\X�'���Y#�� �v�'8����ZQ�Ѱ&AX��|��
��N4�2 YM(<)U�,��< ��7���DōR�� �R��!�ɧ�����T���PHt�����y�,S1���Ju��S�Y��K�.��ת\�rL�@ �o��T$qO��D9E���aT�Qp":H�2ʄ:�!�D�
A���!�L0B
=S ���xe�$��we��p�9���-0c�J����2��DAf���C�I"����R�O#P��̫D!I��F���'i�"���d)'ܘ��M�?6;f��c��	na~��E3a\ip����Z��\'������\ �� ��>��(AT̃+^FX;��̏-w��D|�'� ��I ��BHܧ8���N��xl<�k1�B����!� ��

Byub^= ~��Γ�����d�R"�ӧ���ٺ$옐~�>�P[G�E��"Or�:���u�`�hΉ"�`�ڡ��Ȱ�H�C��0��'������'W0mr�^�t� ��a�,X�͕�<�	�A� ��R@����c8���!�L��
�8U������&=�>?N����� ���>� m�fEڋ=����rL�6t�is5"O������p� Y'+�P��C0�O��3 ��;[Ӭ�O�>�s"B�NP�|�󠕊J�r@`7� �Sb¤����Tḱ>\$	�N���XE:AY�t�TdT:d��ybƄ98n��=s��:�����O������	��b>Ey�H?JNx)�*.1��(#�0D���կ�87��+R�ٲU���;橮>�`�iɘ�څ�<}���7k4fH�Z�������-P!�הO��,I�韗}�jP��Z�t�'�d�X L�2�d��O)��C��b_ h��
�l����'�X%��"��]�Cgq����#�nL�p��F�*���d���(G��vܞtBW���y���(ӧG�}aЬ�֔��N���%z�K/jʂ��5�P��y� ��c�XҠ�5b��@u����ϴ!+7HD���)ҧ�:9 ��s}NtY�m�2��ȓl����3.q�����X�H|�N��)E$�:�ԉ�N|�>��ǀ
>�ZP��K?c�TR���h�'��@�'K�I�P��h!o�{2���!��������R����7�'�l�aO,:�9�$D8����������=��I�frr���N�	��IEf\�y��3�V���̰�@�� ���&ra�i�D� � \�'��ð�����g)���mZ3�p�B��N�
xP$��I�t��V,��:�f��ɘ�=��dfW�k[�ݛLFj������Tj� ��S;tS�ax�N��HO���p�)3l�����4��a?ι[W��c�@@c5��7�~R�=�O��ѡH�6��r&�an0ٵ�i8US�\�_�n�O�O��'Q�I�Ê�c��	5	қE�����'��M+e�#���FB�=�}�'2�8:c��((��|�e���8�n	�C��4ef�A��vX���2Y#h�\M��3*�#c��|�h�ׅ	)��5Gz���'Bȍ�b*�QCN��I�j�@��$ڰ#��x	��(��O�
d�tG�2=ň����b@jɢ�'��	8o�	�5�'!HDa�� Q� ���*�\�r�@��V<�8u�����S�O�F���J�>i�|`�%��_��7�� �����O�� �i�Bh�!į,[�������f��^X�	�tP�w��Y#�Ӻ����E��m��N�)pz<�Ӥr�<��Cu���[�ET#Q$��Q�Tu}�\;*��b!�M���,J@Ђ!D���rc�Ġk	�C�I2+���G@����e._~�,�O� )ǃ�	Z��%>c�x ��D���2`��\��R�2�O�Uʠ зZ��d�0n
���]����1gjNh����?���
�W(�]�q���h C�b�D}�O2\�O�C%Z6Tt�H~BM�;J�@� �-zAAuʊz8�P�E���)�To�7�:����9��x�e�̒Y���>p�Y�R/a�ҧH�b�;�S_�^\�fÔ5C�i��6�8�����Q>I�f��4~���X�2hЄ��
�d��ˍf֮����t�3�	/a(�e�gJ�/L��q��?>Ų�2��؄|l���В>E����Z,{ ��HH�"�"/�@q#w��1E&��gh�qeV5�n)J0�I�T�l1ϓRh}Ao ���':���n�^��]�� O	v��P�qQ�����D��2��.P�.�@��GK�1@��)w&��?D�Dɥ�K+uvPA�$N�&)9��8�$�9�R�HU��|��A�\���B��4	�:`�`��h�<�d"K%��p1F��$���$O"�t�qm�
g�ӧ���31��K�MV�`���B������8�W�Q�D�b�O�S����S<r�!���$�����o�^�I'GN�B)!c���`n�|�Č(����ױi(:���K<-^�8��KKC�|���'[KE�+4�t�w �*Ni��^،Ez"*LR�vYE����
K�2!����x`��<�y2�D�Q�ոW�$^v`qFE+�y"�D0s��*3$��d�*�CN.�yRG�/X�2�kS'_�<Q���yBPc'ZH���I�4�"L��y
� ԻP,�m�|%��G�7}1fd��"OH���iC�7-����W;Z�eP`"O�):�L�1���C��_̄�4"O��'�RĉP:3L��X�"O�"�D��e���j?�D�"O��k"ڱ+Hz%c���3J�0��t"O	�֧SJe@gm�Q|�4�T"O]�w�ڭug��j�Õie�t"O�p� �U�jޠM9��ÓS$�\@�"Oz� f�̕?�RX� �̨!�dU�6"O��aЊ&�f�j��\ /(Dr"O��k�Xʝ�Pȋ�Z��xJS"O����˕�WX�t@��D�޼Z�"O�⒩�3�ԕ�C!�(%���"O� �!�Z�w!b(hO "9Pd��"O"�3� �q/ �J�N\�|� \��"O,�J�k� G��a)W�*�����"On���J	b~Ҙ�Ƀ5I�l�Ӄ"O^� � ͩql����T�:ѶQ�V"O��� N� .��Cu���X���"O�`a��Ò5�\�8%DU�| �H�V"O���6�P7~x�$��0K�9b"O���p-�U� S���1��"O��	+q,��D��#�]�`�	�nL��'C�Oې�A�Ɋ�d�<�1����';��S!�!�؆K�@�(�6,4�)B���"!���2� f��PBj��m�,
!� -ʆ��`��h�Q�
�;�!�ϡ'G�Y0�̃�x���Kh�"O&�)��D�	5��yT*@<Z� ��""O�9��D"|Q�H_��v�{"O�ASa�J�N��	�Cǈ�dY8 �"Od��ç�o2���e�3H��3`"O����*Hb�2�Ć�*���"O�)KA pθ��EmI�:����W"O�<�#���	k���3���˰"O6()�h�Q�ck"�ִb�"OL��Gɹ#���j*C<����"O�Q�A�(_4�Y��3����S"OСhJ8 �d�QB@v���҂"O4!Zq��[���]�U�F(C�"O>����+�|���$��$:�"O������e�I�'H�n�:��"O���ŚNM��!b�MO���`"O���$C�Aֈ��C�22HeI�"O���f�P,M5��₦t.��y�"O��ٶ���䈕ɵ���"!zx��"O��X���=y=^!`�O6.��"O���a������BbI���h�5"O��1!�w�i#a�h:`K�"O��Vꃀ4y&��6@��xऄ�1"O��a�f�!d�{4 B6b�є"O�9��7Dxv�&�
7dkҝHR"OF�٤D�3Ҕ���-�Hj��;w"O�%�q�8w�.|j�.5v�XeK�"O��pLޥ0����'��H:0i�"O���ŉY�QjL|*�� |�:0rp"O���I����eל8�f�;�"OHlx!^o��e���hI	&"O�\���lӄ x&�D�O�ȸ��"Oʍ؂cO�i�H �nϸ~��L��"O��"[(i߂�����>�<���"OF�
D.T�:��5�:9��ȋ"O֨ �ʍ�Ir(ŋW�D2!�H�W"O�  a�� ZG�>8��NN�ua^��"O�e�Q��OH(a�ĉHc��Rb"O\�@UB�j�A��4LZ$Z�"O��
�M� O}�l�V/Q�2.�Tt"O���f�ӵRI��nܫ	�"�"O,�("�Y?�t�qC.k�l$("O���a��G�i4��]�f���"Od�AF7::H3��%4�:"O���e���~o�"3jX�oo���"OX{���C�֠��6d���6"Of�&ւ��i��*��uP<MJ`"O��`p�7Ȍ��c@��$:�9"OB�)��>"�5qW�[�DH�"O>�+�<D?Z���U:T	�$r"Oā{BdE���<7G�\b��"Ot�qR�~�L�Sň�
�297;O0U�G�~X����\�\}��1�j�.��`Ҭ3�O�TI@��~c��D��x���)��y���W�yr�͋z�|����(�$���mH �O�-I`�����@�q�eZ�*l��Q�\��j����:�G�ԋ �J�qB�P2G	h�b`�,�`�4�<�)��<�c���4@p����+�E�0}�`i��d(�g?d�G+E�E��K|dh3��U<b�_�,� �0
��G��qQGEn� ��T
jc�{��'�&��g�׷wH*����.2�1���	?^ �rBПC�:�{��b}sc�m�����@I�t�0"O:U�`��0Hx�d���/Q-��X�ດ͎�&�E2����.��?��1��. ��Z��s7� H,D��hH�2s�$�Bg<1�(�1�L��F��)�'�`�zB喹��ϸ'�Ne�A��} ���EG�.&l��c��U���'d��#���'d���6��;I�y4iįF$P��"�5�j��rW�'S��h@
� �p=��gB�J�;����6͊tɖ�=r6��Y���'E�(p�E����2'�F���T�p�B���dPi�T�V鑸�az��	�0A:]�tX���7$�9Y���3v�(��
�O6?aa��^Ш�
�R1�%;##OP�O�ډJ ޸;�@��_�r�ٌy���[�b���>G��!�#
�.ͨ��S�eU�-�L �%
*G.�ɒj�Q>�bd�;�E��u��<��a
.6�PbƦ@���>�pF��OJ� ��d��!���qôP�U�j?	
�d?�F�F��u�7O@ � ��/1C��=�ƌ���ϫr�j��S'@h��k�*|Q�j��"�tqh�<]t�[�'�@#v�烅�0�p w	�WPR�0j7}B�2b/��1�X�Iw�%6o�˓M�n%31��/
���(5�����$�=�A�Y��l�r#��A\|"<Q�&Ľc��0¥M�(��bU� ,5�B�i4�J(c���f��ay�(� _X)�'�՚^���Ć["	�m�"8rZ���B����U�ԉXu::�R����0O^5�e�,v�,xC�a�0�n���Ec����g�7ʍK[c2,kRfM#��"��:[�7�0�O�3�@�f��:G�I�2�)HҘ1�H?�	�t�-��<Q�%sdش7&�O2A`�ɡ#z�0sc�C��`Y��	�hv���}L�Y딎x����p������ �-�L�q��Q���"�8M�A���DYg�A�˓;����B2z�p �ȣy�����q�d �CG'A�=��ə�{@��>�� N��dl��� ?r��i��îY�!���%�R���D)6M���FAA�t��[ ��0<i&��J����w�nȲD�9z�� �
R�;;���{�����@�ŉ&$;x�q�C�nԄZ����k:1���3�v����h]�i�*t4��S˯=X 9A��i�" 44���Q	ۏ}� 8C�;O��9c��;,Y����f���!�sF��ɂ5Hi�ahb�l�axRH@tv�A���(�Z-��k۫��I	\��X��ǖm
����r� �����^+6�ۥ�	8f�ٰF�O��B��0U|@�򇂽*�e�`$N�d?�Q��4n�(٩��IF�'�2��*ɯ�y�a��Y(�n֬Q��-D�y�'3����k����f�6���`�L�'vm����bV:ECA#݆G��!�O
���ޥLҞ$q��Ӛ&�R�	�'�<K�U�u�0�X�#3���k��P?�d���8|(��3�(;vx�Y&(yЈ!ŏ��s�x�j�<U'��ظ8S���o��'����&/5R,���ԑ ��[|�S�? N��7�I�F�h|Sn��P�!�HH<�ad���p�Ȃ�3V���&,��XƦ	Z�֨hx80a��>}2��U����.B��;srU� @
�<�$]Q"x�Ɠj1@��d߭N&8�AN&Aݔd�O l0�H���(�X�@��lύ�6S I>�d�"���Q�-̲���e�f�az� �6&�ru�6P;��D΂����Fo�-Jv�2Cfےad,��Dhۻ-t6�p�l�s���$��"��㔆B���ЈD�[�Q�H�%��f$�ᐎR�_!�ъ@��OҨ)�"��{ \|u������Ʀ�	�ē"}�}0�EE8&7v���	}��n�OJC�֎ 8�4@0�ߴ��7�6Ua��)�\c�R8��bN�R/�9�*)�V�h�'|�y1$����J�kF(-��kŔ7��x5,8�ɴ���K��z\1FaQ����l82|��O�rښd�w(�=���dN	Ype�L;�H���@:>�b�	�J�צ� �i+; �J�D�~A^(��6�f���A�ڵ�
^�z��5`�Ù�џ�i��
8�� �ӈUܟ�@���tBBl��<�H��a��/����C�dD������m���g�_8N
�M����Q����k5}Ri�V#@h��M�ʟ�	�A���D�k2F��c��qߔp������L���B�$i�E�K:�~�Z4�B0��۽U��\i��Ҍ{Ψ�A��Y����<�g�K3pMB1�ORQ�u7�.ak� ^Ǫ�*b�M�@�.��"OD4;WM�)5�0�q-ϲN�����OT�3]����+��)��J�%���Éo�d�A]+|�����b
�U�6A(�-/�O�e�I0f�zm̊����O�,�牋wQƭj���,OyT(¶		$Z�f#>)e&A��0���ӤT	��C�C�'�2�� ��&R$��G.�J�K�
�t��A1��^���])��  '��KB
4CKa~�	U��0�"JI�QpD���E3��d�e�F�u�ΞVM ��DJŌq�S��f��XB��HA QH������6�yFq�$%��Ŭy����:8����BB2�\ͤO�Os<�o��5���7����oO��IB��R���R�=w n=���:L�B�cq��.-�.0+�1OZ��`"�V�h�ж��"�n<��ɰ,s��;A���q r 	WB\�?����z�>Yy�	ءL�\s1$�<,}��HWo��4$Z���^��y����4uv�J�b4�x���Yt(�0�E=�$��'�dУ��,W��ّĪ��x:N��'�ƸJ���?b��{��X(Z\�ńȓ3h�b!@�F�0	t��)Aɺ��4�V�dk �sy��)��'$��'@�zbMTGR8I�%y��S�'�\<{�̘md��Q��'�,����і�΍�BNY;%� Q���%t�B�B�?J��Ec�dBW�P���+e~(����I�\@@�'�s�m&{"� F�ԍI��'SZ����N84�XY%�x���@L�೶B>q҄˅`Z+W?u���ʮk�����bԹ �m���#D�\ @��"( 5�&(M���ݓd��%@$`+�
�>y�����'����K�BNl�D��XG� �'p`� bW�~�P����(:� �[�';��i�����=�Ң��`���.od�����s8��G��;L��m�

��lX%nB 4��P�������D݆`A��T_~���\�>`��5!V���o��O��b7Z!Q9آ}bB��E�`S�+�40�5{���K�I�mp�+v�Z!�0|�b�)l&,%3vBװHi�hg!�= �6��b�B��S��yREӾ,���F�YNd���̩%]$͋J<�SțWC���'wfV.L<d���K����m��'�� ���Nb؞8P���[��(���� *8<j��2Q�lQ�����p<����vy�_�x�&�Ҧ��=LI�4�'aV=��<�&��?HA��O:�2b`G?�\��!�@�-�Fd� �'3��!eb$���z����O\Z����.�jC�	�?pD ��Eƀ+�-� �T�D�_0�;�)�'U/$,9�`�3ƽ9u��m.C��;�J��w�O�'�p�r��g��b��2���c��x¡��܎���̬\�����Ù�xB���nLpi�J� ^"(�4�K-)��T�g�U(<A�Hb��bA^#l���@N�x8����?��'���YsH:(q���p��[Vf�0�'�9)�k�G�25���Um2�I�'�L�4	��-;�|A�[2p�'�$��@ۂ]��_VYBPS��� ^-���i˶�"6,�	^�6X��"Oew�E�|�<�WKW�V��ja"Ovă�쉜x�p`YV*:����!"OR����	� $��/�^p��"O���ࣔ/�i�S��j1ht8"O2�YFAZyeB��L��g0�\�"O,=�!��;n$4�k!w,��i�"O�h��SdY��T�=Bm��"O�YY�c��ZKp5H�Φ&<��"O�Jr
��h��N;=(ũ�"OV]�ӌ־S�:RG��Y$��)�"O�8��ȂL��ͺԤX=h��"O<���mݶ'N� �ۖk2	�"O�)��N>s�DH��S%d�\�#"OU��M���<My� O�?��ѐv"O��"LU/9�4������Z�X�C"O&l����_����Z�����"O���Aϓ�	�8����E7[�n�z�"O��2��L�ص � �3Ot�@�"O�|�7���K��$x��uj6���"O����)0U0�b�O��c�6��"O6X:�!ް �MX��%�� �"O�i�O^� ��d[Ad�1[�QS	�'g�=����@J�
WN �R�P	�' �Z�D,`�8�	0$�+;w|��	�'�<��d�*\ztl�r:"B�c	�'�|�SL��z�?#q�I��'^�[cBӓ-��)Ys�J�>a��'�.i����=h𠋢��7Ј��'+xt �ŗ,Dhq{A
M3� ��k�h(Y�� ��|�Iܾ^Ȇ���Z�E��A˗u�f(P�'�Z$�ȓ7E���K]9d�Z�"(-RFa��O�`��G#�%&I�)B��+7�H�ȓ �� Xd�(B�fJ��8\h�ȓR-�1*P�H�d;}�� Z�%G�'��z�k��p�*ר��
P���	�'��M���X�f����6+��k�֠�
�'j(���d�~���tn�`CČ��'��&"�D�v��e�֙P4�8�'T�����	�j�RUK�`1�'��� 1	�[t��J.��i�'S,����r�r!�̓�G�t��'q�ר��+�N�`��*6x�s�'�v�rf�J.#�Y٧�Ўu���9
�'n�8;��,�~��d̏�6��@�	�'�@x�M�,\���%�& ��a+
�'�PQ�ƥӕ/���{��vf�q(
�'ɞ���H���S��
og,��	�'{��p!�ߋs�H1�I�f���	�'�\��U���н���ΕZ��j	�'R��k$,t>����O��i

�'�@��O�+H�I�e�E˲�	�'���J�c�$: ���'�@44y��'d����!ץ_��  @ު9�d���'L@����:f��<� MԽA~�q��'�(p��,�5ot����/�,�|�
�'�N�Q�eU'%n���g^�j�"	�'m�Ѥ�?��%sG��D��S�'�f�r�X�87f����̚h
7"O��p"�P4J���E���3ҢP�<!S(�GXr�+%jݼI!w�_W�<!�K�R�b�C+�v(��0�Xm�<�0$��	��MT��(1��&Ol�<� L�!`�Y%3��9@��:^�8��"O����d�#̠A0�̄R�9�"O��8fB�0��Kg▌I\�q�"On8�,�)!ϮE#��{���"O��.߯N�xԒC�K�l�&U2W"O�䒓�N�Z P�J�(��0y�"O"|�v�[#R\��CIA9mt. �w"O�$���Z<d �
(W�B!��"ORT�ʊ3Qv� 	Ӈ�:LVa�C"O�9�� B"rЗg͊yU̝ɒ"O�R$�?�"���L�t���6"O��Bl։5K��(�:?�a�"O>�ӣ@60� w�"�U"O�đ�(�	,d����O-084��"O��2���j8;� �� ��"OΙ[�l�4=b8������Ib"O"-h@�@�~�P��ɄX�H�"Or���'�h���*١MA���2"O,`��J�2x��(-}$XЋ�"OB�:t-)f�.�9E��$j8a�"Oj �NP.jD&R��X%'��\qw"O�	J���'/�d\� �N�F|ز"O�LIq�|~X!q
�!˜���"Oz� �5D��۳Ӆs��""On�!�k*@d���/���7"OF(�C��9r��Cր�]BN͉"Op�Yqb�?i�T��F�VN3.E�r"O�X�P���8>�� �@8/�y��"O��I���D
zQw���5��pФ"ON�
�#H�8�V���U�l����"O�����0h��!�BW�6d@2"O�t�G�]���AG,S����"O6Ļ���@���nG L�Zd�d"O�)C�D��,�tZf�o��:a"O�<RVh
+J����K�_܈�.\H<� ��&����!�B(D�����@�u؞P�=��K�8W�a�!�>k�p���M�<d �@�h��F�ȗ�X`rAOI�<Q ��'!��@KOȻQ�u�wɘB�<ysH(�J�"g=^����~�<����Ѐ�e��%i&�C�a�A�<YG�Q!��e�J�$e�=f+N@�<� �7W��p0vIc�h���~�<�r+S`}�t$�ER�x6C�~�<1RL��P\��:t	�,Bf8;� O~�<�ׁ�@8BM�ċ'
������B�<Q'�͑>���O.@aS�A��<9AI�/G�(!rt��
�8�@ʓ�<�3�a{`�EA�i��P�oAr�<�t����Ѫ��(h����w�<Q-ϙi�����7}��#Xw�<i 'Y�QD�R�W�|�2|�è�v�<�r$���A9!�L�+JIxUs�<Av�!_�(��ѕ"Q�����e�<��A8!$�{�Oy��i�fFU�<�G��U��Ԩ��T����d P�<i��l��f4:5 d��ȆB�<)�,�E0��d.�5b��T̉�<�1�T�1$�ň�
��!j=(#g��<�AE�'6�C��Ӗ@�d�]}�<y�bI?kXȉ�+�6_���dW|�<��R�23N��`[�V4vls��t�<Y�햸4>��ZDfV>6�0��o�<qqj%��2��=Oô I��h�<� `����3*�`�n��\G�$�"O�0*��W"�ʣ(Ţ3�hY�"O��2䨗9�:�xq�Z���"O�Tb�H�K�D1y�E�9h�p �D"O���%J�����YcD��S��ʕ"O�N�06�ޘ�d��{��C5"OzT�s59̀	CKǅR���#`"O�D;�DJ$✕"�i�U��R"O��G��+��Y�sh�0k��i�"O�M #a»M�Lp���N��!J�"O��@��%Pl䚠n]��8M�"OF4�A��<��q�umKj�j�� "O=�T�2lm�����`5"O�U9�M�@�\�۵�LbS,� "O
Չ�iߑ
K�����2K~�s�"OZu��H����� �gE&-B��
U"O2���&.�y�ą�[AZ��"Oj��G#�SE�Y�RB��@b!�"O����:O4����W>^x*U"O(�pgwF�qP��?6�0��e"O��P'	ܣk�j��w/�"'���D*Of�����3�D	���I�H)��Y	�'1�u��@0�0����.&����'��:���+r���(�"E���t9�' ȵ��
	S��p����}k���
�'Qҥ#�C ��h���6wU<�@
�'��5*1��HD0r���xN,-��'�H�5��;-^X�C�"v�B���'l���v�B)}(�����Y�)p	�'?*�JW�A� 
~ɈV"�!��	�'Kt�ZԠ-�R�+������'6�=I��C7 �&l��Z1�
�'��9�5![�ze����v0�	�'�����΅�W�R\�$M�������'vd f�кb�\�"�� #a$x��'h��%�ݏ'�إ��ϕ����Y�'@X�B�)\,�RǛ�@M��'��q`̗1R1�	��M�`L�P��'5���� \Z*��H2fL�]����'�,���k�)Sk:]X�a�FE*I��'¢Ԣ#�܈l �C�/�A�����'�PT𰤊5���p���6@8��'�*�qRC
��Lي�^8����T�<1�M�468��-<46t�(7BX�<94�P�I�J�GNGt{wd�m�<Q1�ԩcOt���CJ���*��l�<�U�Q�k�R����5s^0�'2O�RD����� ٘m��Q"O�p� "��p'05��oҸg�*`�"O�P��h��c���SO��h�Hj�"OF��3��:Q >ȑ�m.�XȠ�"OB�AA��TY���V/���8r�"O����kF�&X5�u�:�n�q�"O8��!+�4����"@�b"O��Q��*H%�BO�|� "Oy�&���@c��FEƅq�4"""O�(�)�1.d��Ed)9�䑇"Ol��u��<��@ !�ԫd� ��"O|k�+K� (��3T�I�O�V0(E"O^\��-�!S���AW��>���"O��w��-)��5�&/�/�8\˅"O���aBU�D~
�r�M�9*�|�j�"O6SI��.��KH�;�d��"O��Å��5����'$"
|��"O� �%��
�(1��%E5x�8И�"O�	���_K�0�
�MFb�z�"O�P�c��OU��ʖ�X4UW�+G"O&�����?3�ı���f>2}�"O��#���l-�|�`K��ON��3�"O��!bB���1���ׅ�y�lG��q8gn��z�|��U��0�yҁ�%L��A�p��@!DmC�yB�� ��y��o��j.�	���yr�W��1ӪY�e:(܃��,�y��ˣPf@�ug؏YǜL�u/��y��v��`��Ç�e�h���@=�y�W�N�� �A?c�Y�ǥB)�y�
;.�����NP�X	�����2�y�����]���.hǮt2 ���y"!�g�+v
��Ys��7���yҊ(kv2�ӅW4P�8��֥��y��9}cGu� ������y2���%����H1p�$C$�-�y�(�;.y|XA_a`����ח�yRE�XQ\�ǣ۔	��iW$ (�y"��edq��б~%
a ��Õ�yba� M�(Q��
�v�C����yR��kj�Y��B6~H��qh��y2�S)�E+E�4-�:|� ڴ�y��&`.$I��B���9bvkP��y�7Ob�i4hΔ��`x����y�b.��޶\8��TK��y��͹c� "we΀^3�];$�C��y%	�x3$H���/^�Fq�0nT��y� ���L��Q�V`�{Q����y2E�}������3^��dx��H��y��F�Z��bGM���#�����y�#�ot����2麨bD�^�y��#c�peÄ��.�{�@(�y�H�&,nr\(���*��
֪���y�'�,~� �imfX�eN���y��КY�\��f�0>�b^IV�B�ɪ7��=�S��#uOJw&�=)��C䉧`���)��^"du��/vc�C�/0�xP;��Έ0����tA��B��C�I�5&���-Z�A�c
H?�C�	h�<�g��W#�ْ�*62�bB�I64ؕ���	�������orB䉋]�h���Bŧ:纨`ԫT1xnB�Iw{��O:J����Q�Q�DB�	�[x��4�P�x!^$y��,Y�B�.� ��hAj��U�!τ%��B�	m`~��w.H�j��yh�*�=�DC�I8Y_\��f���D���)ño�fB�I�@�IEB��W�=Y�2> JB�ɴq���Ye�8SI5�Q�R�]$6B�I7 ���#��NN��z��>��B䉞����U}沠� �N:��B�#Sq6��&,�H�D��g� �?�B�	s�t����mb(U�B ���B�I2ZS�p��l��4����܇+GrB��3������ "��ر�[�`f~C�	5ڹ��͝#ʀ4� D��DJC䉘1��$�3��Z��H��4C䉪Fj��B�-nnq��!7h$C�I�7%($3P��th�R�iG�	�C�ɿn����s�1��UҴ��%C!2C�I�8퐁	4���	F�]HэP�:�(C�)� Hݐ� ���t�U슽jr�k�"O8� ��J?�гFME���T"O̝�Q$S>BL��W��IkZ�2b"O$�˳C�ބ��1DU�)��"O��¢ꀚ+�0��*�:��9;�"O�1�T�%B��,��u�d"4"O�4s��Պ&���a�
����"O�a#�U�V�Q'P9~VNu�"��XG{����PQ�Ȣ'o��ŀ���� =�!�D��fn�V	Q*�4���/�!�D%� %j�c7	��H��gQ]�!�D��I��`�"�=o�80���,!򄍐\���Af(D����6e֌_!�Ds?�QCC�ClfµC8V�!�D�|,�T)C K���`xS"R#U�!�ݍ,~���,�}�Y�G�-|�!�D�@��P�˂a��9jEG�#{�!���?�&}  oψN2�9iA���g�!��� o��ՆT,���Dϟ>!�DȔ]���3M^0_

Ԥ�9�ўT�ᓫ&9]����=DX�0��,M�ww�B�		L�e0Q��f|��FFL�:~�C�	��`d�Q�fNȑ����B�I�<�qBQ���c�,�6j�H�C�ɀq>�dH�|**�ґ�>v��=	ç;����\�-�p�@�͠[��%�ȓZ7,]�7b6_��4�w��E�؆�n��H 2�#��qbr�D�BB�ȓP��T���̳h����%F������������b2�5Y@��m'~a�ȓ+�޽�2k�j\i��+�"F65��y�����芼L�5y%�L!�2��)~囂BED�l��BA���P����K��^F�a����"~����ȓ%�5�	Bg.@X5�ɦ+�J��ȓ%T�P��\�ɓ���V{X�ȓ��y� �6	(b���]��ԅ�\~�g�G�d��q�EhX�!"Hm���j�i���RTò`N�	n��ȓ]�.Tc�	ɛwfҁ����K��ȓ��(jc��$!� �dݔ�ȓ	��5�� ų*�,�1D��(��ȓgtDU"\-I�z/��% Zq�<i�N�1c��q�m�-&�JB/�n�<���I�v$���AΦ���%J�k�<	�+��,�����ʟc���7��f�<t�P����1i�hӸ�B�	n�<�`�� Ą�`S��+W� x�5�CP�<qs��p���3�Q�D�ɤ#w�<� ��q�"�V��1F0����%p�<	��>ny�G�܄|\(!�ˇn�<��ЂRex�q�MɬC!p|�RD�g�<�J
]qJ��QO	0!⸅�b�M�<i�l@)0���IeF':�b��Ja�<ip�?J!���f��=|�[���Z�<�e%Sf}T���#U�b-ӳ#Vp�<���	0���6	�I���·��C�<��N�W.�X�Ǖ1<Rs[�<	����*��MW}0*���g�~�<�5 J�9�T�*�"%A�<�gT�<���{�n�x�<y�|�m�R�<YA#�FcX`��BȤ����NN�<1�a�
��"3
ԟd�� (va�I�<!PO�M-F���t��{�`D�<� ���7I�����c��4N=�<i%"O��j!��2g�#o��`6~��2"Ot�sU�<h�|�PΒ8*w�`��"O��ywL�J����W�ye���7"O��H���E��{�-�>$M�I`"O6=bUH���hP����+OءZS"O�(����7�*D+�͛/#H���"O�	i&��}�F,KRU
�K�"OĵJ�B%u1�����;C���'"O"�ɠ�B�H`��̆�CN\̒�"O2e��-
�T�!�3lL�?�t�!"O"��f�V�iP�+ .
��g*OF5F'X�Or�(� ��;�'�tAR"�ӅB��4�qF��
���'�)�� kd%��IFs�:0�'MhJ�+�7S���jumۀ`��s	�'2�tЯ�2a�̈�b(TM���'&�4ڧȏ�6��H��U:� Q��'�еY3��gG �KQ%	�2Q�!��'7V�#d,}�^TϞ� �r��'��k�N�$+t��肮�^1��'SP��Q�H/0���.܄zH���'���2�Lw@~�%i��y�'� ��t��d�˗
{���'�ЅP�O�Cs����>	&2��'�������'�8	q�ݼ "��0�'�rDC�NʓoԔ͒�A�&��	C�'����E%�Ph��8h+�'�P�k� ��*�D}P�������'�\a+f�m  �kŽx��*�'�r�#u�<�ڄ�2Λ%�&̓�'������
E9��I�� r>8��'$�t�@m�8���+�.}�����'�*,Z���53��B�/�}b�`����Ў N�! �́@ft�V@�)S�!��3b����G��,PrҮ�(&�!�DI��
D����ֹ��/�:@�!��_�F(ݐ�BM�I�PpHF�߼3�!���	I�	�R��H���J�!*!�$י,�j��HЌN�|�3 �=`!��Z4iA�e)��y��T���¯!�d^�4]$�K���3Px��8�'�O�!��(%��3�9Ddn 账� �!��G�q��h��JK�f����K�!�d� %RK �՞{�PpZ���6�!���F��%
Ga��t�(0�Ԣ�?l!�L6$�D��p��x�� ���C�&e!�$˥ʀQT�s���P�� 8d!��=(=tL��K��O�"��L;5!�I�"����FЁc6���	u!򄘪|�L(+��-*;R�+��;ng!�$�0@�B�s��Z�A5(�,̿O!�DM�Z���P��e$6dC��E�v��zr�ibBO,e�Ui �DA��O="��xh"O&���d�%x�MPg�E�\�ɒ�x�IQ�wɪ��V�|���$V)p��=Ү�u�P)���y�L.���#�ה�`U!̵b qO�`� Wq�g�I.f>R�ƠG�d����׃.��C�ɧ6-��DNB
OD*�2�I0z�~C�	�-�z��ӦS3qD0s�Er{�C�ɮ9:R�M��d\aLC4����8��T�T�QAd��@+�Xz͆ȓ�ƴ�7�ц8��b'ũ�� �ȓx�9
7���DҪ�3I�������S�? ��e�O5bk`��u�\�/���h�"O��"P~ q���3w}���"O�l��\�3�RP��&ŒD��"O�����g`D�7��=o��e�C"O� ���:\��Њ��?���6"O@�k�)^hx�Q'�
�6�{@"O
�rj�I��
�FR�"�b�٥"O��h��M&nF�q��+���4l��"O�T�+{!c(_�w�B�@�3i�!�DV��� ���v���^#�!�_�b��rs�������`��T�!�d� a�F���P�{�P�A��	��!�	R������SF��Q�#��6ka!�DX#8<h��g�M�/��P#1�@�!t!�D��H$��ɚiN����^�O;!�Ŋ}5�I{3
�1b%(WI��!���:>�
E��;)�e�g�g�!�d�ˊ8#v��27��c�n��!��J,K�}�f*ڥ6�DY����|�!��10����EaT�J�&�P��Y�!�Da���ѦS&H�`8�qJJ��!�ę/pV�tr����b��̲DCѓ|�!��z�0|;0ӭBQQ�+e�!�dtȌ��w����$�d���Py���am�����0#�K�hF�y��ƨ/zH	��+���B��"�y�Ч��a�aD:TA�J��yb�ϵ֪dbf�͕NF������y�&�"-�z��ŭ�>1��mն�yb�A�.�����ĝ	����ҳ�yBɂ ��S���y��1���y"-�+;��p�D*�v~�����y��M�D����-j��0�A�M�<�s���Gr�4Z�@�1
�Zb���P�<�6`��m��BN�1'e�]KBm�c�<ѕ�T�s0���)�1�TK#��w�<1�`�W`V��V��Qo�0���q�<�c(ǛZ ��)C9|ܔpQ��h�<yrG�U8v���	�m��'�NI�<��@��[*zirF��/�8�ʋK�<1"C [�`�c6��4faS0cc�<Ap��2�,Q�CӅqoV(RmYX�<q���1(�)ኛ�a�J�O�W�<���\k���b��:^�*r�U�<��iD� ��� 6N��uB�Kg�<���Z���Ѡ�
���="�@[�<�LI�Mʊ�I�G�h����nC�<� %�fg�(g��d���1�CJt�<�c�
�+���@�̍/�a�p�<�v���,�&���[�H�Z(���E�<��lң_���Z-p@ҙ�Q�	f�<Y5e��}�A��c^���[�<頀�5wm���FV�>�Ex��W�<���
�w���pq�c� 6fU�<Y���/0�ި�b���=(�(���v�<�cOQ1�l�2!L���q��)T�;���%WXȽa" i���R��5D������u��@ZF�C+1����"*O���"��.��8����BZ� ��"O6�K�F�	�(hYe��nh��ӳ"O�T�!�C!9�#B�[�Z`�"O���Z�$%Z�-�U"O�����9[1�@�^r���"Oz�vGR���u�M�6[�>Hj�"O� �H��h:tΤ��ŋ�A@�a�b"O~�[A�]&M8��k�;J%��J�"Of\��ɗ��)I��S0}�({�"O���#Jф!���f�l�v���"O��h�lI�#�& K�N�#F`P�h�"O�����̈́`��AS7��P[��B�"OteaP���K �`�J�SiB]�#"Oր;f������LJ�i��8�"O,yzC��T�t��*��P���"O����Υi �|Q��πzM�=J#"O<X����}��Q����h�x;�"Ol<��c�6!�zR�]/��A"O(��1��e`Z�s�NF�AfBQ�"Of�E�[�Av�5�b�ıKF0�"f"Od,��CY�`J�Xʆ��46R��"O�8A�`������eU�]�"O��� fQ�,m�a���rʱ�"O�$x'�܃�R��f�I+%�D��"O�<�Fa�4���)�d�S� 1�"O*���Ù,v\���D���%�*��`"O�x��A!zD�!ۅ�C9�~4�F"O �0��0��i[u��-Z����E"O�z��W��0�zBA%Mx��`q"O��P-B�i��@�b�ݬe��"O�pЀ��j;܌��jK1yHU2"O��#cC�g;�51��T�!K��I@"OJ�r��[�W��i�6��`:�Z�"O.<Qw-D�|�@E�)�s�"O�TA�́�G\�a��J
-$�1��"O�<Q�%~�����H]�	
��	�"O�Q���l��K7���|�9�"O��A�D�{�u[&�2}C&���"O2X�l�0\���֡��2�U�"O�p�f	4G�V���c�+F5!�d�&�<�
��B�Nd� ���-~!�D� ?x|9��k\�|#�1�&E9n!�$^�v-H�[�D"�	��DK	!�D7�|��Ѓ��b��Q�GDY^!��R=^i�d�`&jE��BߖLB!����%�� Ł'J|i"��8m!�� L�))�'��+���3F`�	�!�]�a{|����#�8���\��!�$�)����π����1`��p�!�Q�v����Ŝ�"�Z����Uu!�Z�M˶����0*O� �[!��K:1��r#��sfI�dGס+@!���$F8�d�Z��y �Z�
5!��X� ;�@��u���
+!�$U�)E6O@u0�ŉ��@B��7Y�����$�#���2�S� rC䉤-]Ҵ \�9�ѫ3#ӵUvFC�I.Y[Fd����;���K�N�b�C��!i�i!�0 �]�ꌺn��B�<�mp�(M�z�l�a���p�B��G�9w�,"x$Mɳ0�bC�(��u t�ا_�tx�j��l^C�	�d{��pn�#\L���=<C�I	c(�]�F��_
�Q(N̜C/C�%���b�ӹU�c�Ȉ�Z=�B�IC�|�9��� �I"D�ǵ7��B䉬J-�e��*�!���h�aҦB�	�O��[� �r̪A��(6TB�i�p���=8SӁ`�"�"O ,�&�N�.y�"LS�d��]�e"O� <LPbID�l�b�T�f~
��"O6{�@G�J��Ij���<4�(-c�"O$��D���`�I��
�t�r"Of<(B��2Ҿ���!M��t�"O2�q7���mx� ��8%?n՛V"O^�b2�W�__x��'�V$t:>i�"O2���C��22�΁uX���"O4P5��j�<!Df[�b��d"O��U/]��J���v!*�"O�i
#��Z�`�J$��0s�5:�"O�$;@�āeN����T.u�X=C�"O^t��"[	.6���l�D��2"O�i���(Z0�i��J��A 	�"O%ɵ��ü1�g/-h��U"O���1y��
�$?z]���"O�10��̀r v�S兘<dI�Hr"O�.��w��d���/?X�s2"O�i:���B`�So�?T70��a"O֥" %E�o�89��,F'��X"O$��4H�[
~X;��Ǎ9y.A!�"O�,����3-���Q�i�%�"O��ض�J4���G&��"Ol$X�V�g�%㇟�p���"O>�D��d�:qÀ샯5���
�"O�<��P��<��Ḱ�4]y�"O(p���ǃ�����VL�6��"O��r�'��$rV)�${�<ȗ"O>�b��R.>���iB��b�l �"O�,H1�vȱ���n���p��D{��i�,s
Y�@@Q lo�$P2���!�D.;~|�p���Aq�!s����!�d[?,���¡t_��S�-���!�$R�/m�4Y��op\9��	#Eb!�d��W��h�#CLd@���(ڦ_N!�M���)%�ɵb5\[3h�"c2!���(ݘ(,��u����Ú>2!�D�@~��f�T"���P�40!��īa�ʴ��$�L$�u+L#~!�䔊u��={4l9[�<�d��or�8�O��"�N	ۮaBc�Ի�Ra	c"ODݪS	�-0�z���4e3"O`���� �z`�)Q�	)�2��"O�d1 ��>e�L�k��z"L��5�'�'٠��)H�E�$T(��qK�'��&�
�T�4�zag�/R`��y��)�S0_�n�yi�h�Tԡ�M���B�	!FeB�uK�.j���B��	�Pr�B�	{�D�& ���I �B��@g�8s��=Ag�m�0�B�@x"C�əu�Hԓ5D7eШ-�Ө H��x��'��O>�JÆBUP�!-S:n��e��4O��=E�thFe;D��+�}�!����ķ<�I>E��P/�$劁�k@\��f���y����)�$�
�%� �yr�ݔ0¨PsR�-�ƐJ�.�8�yr���+���'Ƕ��%�S���yBI�-��y��
���k�X8�yr�^���y�T �)8d��&F)D�r�|�����+AvrT���)v���WD�#Q�b�`E{������SȬ:A�:v��T�w���y��(s����2%t�ژ�C��y���?zո�ҭ5 <Ӫ�-�y�R�CؔJ'��	d2����:�yb�J�-s��KG�c��a�՜�y
� 4�*��r�т�AS��5!�"O��*�H�{hL�G`�>��$�U"O~�P�:"<N���(͗c�z"O� SQ�J:8�L��FA)Z��I�"Ocp�^�R.�	2H�;8���v"O��AF�>&Ȯ�2Fd��Zq��BA"O8����ѱ�$����cvX;�"O(��C*�sE����B��4	��X""Oh�`��l>����l�� �"Ov��n��8�bh�e޴��2"O�	J� �0p��N�+�\:�"O�a����H�X�Ċ��S�n ��"O�xgע:>ZѨ©	�h�����"O��� ���`d���@��8~x�B"Op\��F\L�!aC�G)`�,�"O8�2��V��u�$i�27��!2"Oh�b�k�����E�)@�I��"O>��`�˔d�4���JW��Z�"O�2�<v)^E�ԭ�6&Q�iB�"O���cG1qI�M��Q��ڲ"O�[�D-Xhx�Ħy����'1OJt)P޵����V�S2�t��'�`��e腬zpM)FJG�Q.L���'�rj��tTD�
֊݂J4$���'I�����n����H�ĩ��'�nHC�± R�1�O�1�d��'xX�����8i�@$"AM`U�c�'|fʆ"�et�􋡨T�Xpԅa�'�Hm�AT��R�ZA���H�:q�'����pX�	�7FO(C��q�	�'FFI8��W:4j�3�d$<�Ό[�'�hYC��������7�*�y�'V��BnM!��,7"P#����'l�tb�e�D�hic���7s��\2�'%$�2jR;�{�(^3oXM�	�'x�0�Z�,,d9���Y�X��	�'),�Ar/�%@��Ao؞%�b���'�4R���4��B��)�h�+�'�b�Ʉ�ǷBEb�J_"�bL��'�<��5��*}M���L�0.BT��'�9p�D��[.ve�L���F���'.�!`&�G�4�K�� _�21��'dB����6m�K\^U^��
�'D���}���*��]��}A
�'��q�Ơ׿S�!���:���	�'��4VKY�>��R�Lh3��"�'���ȱo4
��G�d����'R|�j�,[
4pպ��̨b`�ͨ�'���d!ϯXWvTV%b�E��'�bc-]�q�bY��6R�.b
�'L�tSc"��^�ԓ��1Hb�p
�'��c�-���@����O��$ʖm$�i�q�$X}v=��\?P!򄓴t����g�<ɮ�2'�(!�d��n)�$�c'�)�x�Z���4!�d�z�Q,M+)��Z�$\�B�!�ɴhl����[v�h��I<{Y!��_#%
Ƶ9��ag�ܠ�䟑O!�݅B�!�E�([n&� �A8!�d�]!�n��cR
�c�&!���B��|Q4"
0��5blV�y!��l�(en%2"9�jF5�!���c�$���ႀ5�� �Jӷ~�!�E�S6�u5��:bw�Y��m!�� �q��!X��aV&�x�B`Zu"O�Dx$#Q�&N��/۷�>��"OfqK�I��XZX�Ս��M��4��"O�-:���
	S<� v�&-:1X@"O��q��]4��2��^.v�j�:"O�M����U�ɢ�"ӦH�#"O��b!�ú@8@ШP)��0N-�P"O��J� �A$�3viYx��A�"O�u���$�P{�$	������^�O]L-�d �����I�0`�J���'�� �C�߷Pj6�XF��Z�T���',0$�B��-^ܳU��>�:��'s*u���]�`���Zք�^P�� �'�}��d4d�"��؜~�zd�'<՛�螡.;�!aŠC�|&��O\�=i�BCD&<*@9G��8dj��̴�y��� K㦝0%�|�F�4�y�l�''�]�k�� �(��
3�y���58�I�UN�0�2I�6A�1�y�fX-tT�e����)\�C�_'�y�bEMVL���D�o��9"���y��OHĪ�e�23�W��y����>_L��pm�3Y��D�"��y�cK�&�LI�4�?'�)��CV#�y��	�"�B��#l��<��(���\(�y�b�%R�ne2�i�c@�u�7���y�@�$�}b�O[N��%�sj��y�KG�n���0�U>�8BS���yb#�z��{&�0M<�0�y�F9<PN�:9z�(á���yRiM�`m;������aY�J
=�y�e��]
lm	TCX�J��9�y��J�l���M]�>diXB,��y�j[�l,�l{s��;Z�`{�h.�y���c֜���
X�@�$�q�O��y�E;t�pVË�14%s%aK��y2A��t$I��DY03(�a�.I��y�CB
.[ZɉI�>@���ǁа:$���P�.4�Ijc�+Y� 	^!�ۯli�Zo�tW5Yq�G,B!� �@qSBg�NI�#T��&;>!���61���]9�Iq���!���b�7�ִ� R>�R|P0�'h�ɩW´��M�����fF)V������������<��p�^4?()E��`h<yH�H�$+��:D��R0�OP�<�eGK�:f�<{UC8p�.�b6M�R�<�`�Ǩ|Qt��Z� �bF�D��ȓ!� X!�i��u+��{Ą�S�RA�ȓ?9HM9umPo�͛�M1b�(؄���?1��ڸHᐨ#f�o���7	CK�<y Ό�1Ԧ����D>i��H��E���x�^�Q+2�ҳl� p	�,�&��yBK�>֔�qq�Z=�H](Bd̋�y"a"u����Sd2.����c���y�ݲ!F�I`� �6�B>�!�d�=W����deӰs0�PCs��/g!��dU����/�O��P1OT�=�|���5x?��	��Ր0Ct]���h�<94j��Y��6�
8߶d9RgRZ�<	�� 8�ᕫ����R�'U�<�PQ�����fR��"o�H�<�7Hߦ���)�鑆����D�<��,ս+��Y�rE`üԓ��LA�<� R�yvoɊ>���sA �o�,pb�"Oj�e�E8%2JB�N��n��|j��6�d�O����	i<r��dKL�L�4\y�c�#�!�Obs��R�JYPy*����!�dǂp~�=3�BO�$`���ǀZ!�$��~�fi��ѯݴ�@�$x�!�d���Դ�&���'+D��p#�3 !��]�g�
�f�c�tX v��E�!�~�|��E�>��l 5a96��O��S�g�o�v� �P�Dd"�==��l�ȓuz� B�㒇l��Rr��I�"��ȓ0G�4��LԬ�P5SE,J/�d��1���A�I+9xk�ߨA�V��^"h��3�X�pH�Y��V��܄�.�F��$��-����O��<Ȅ�	Yy��ǁm:�@��
\�*�	�C��;3�'�2���Ϙ'-�e�Kk�,m��ñ5�"`��'s⸡�c��/��� hF))^j� �'���`�A}���KP)�$Wk�]k�'s@܀��_�M�Ԛw���Q	�'��� ��Ѳ7<�QǬ�)���z�'!�x+5Y~����a��}�Z����d=�d�O����A��C|l �,[�G�,�@%"O�1� dԳC)��B�J8 K�ܚ�"O�āǆ�2=2�Q����OZ~�Xa"O��Qf���H'M�:)=&�(�"O�u�E-�8j�	�r�ę%z�!"O*� W�O�[���ŋ��9��)�"OY��eF�F
���E�G�	��vy����_}6ܡFl�^{V��E-PO!�d�/[ >d+��3wI��¥L�%6!��{�ࡱ��͖+����
�a!��M�̔y����k���!1��!�!�$�68H�t&�(7lb6/���!���$^���ˎH_p1ۇΚ+!�D�U:#�$M0Dru䍮B1O�ʓ��B!�੒T�@� �#ۯ)[�!��"O�3��#r�,`A"]�<7zѳ�"O���$IӪy˼��� [�&��V"O���$DW<X�f�
i$r�h�v"O�h���&X&��G�s�+s"O�)
�$`������s3LT*�"Ord*�V;A��a�����c"O؅�!I�?t�֭B���<�Za$"O~�(@��|J�C�ގ�ր��"OV��^�OM���'��}&H@"Ou@0��9ߖYS��>-��@� "O�h��M��	��S�z���"O�@�IX�Z�$���/h�0	k"O�+�a*w?\x�cѬ(�6���'��!��%�˿t(�	�mîa@C�I Y�ѓ/�Z	�4���A�Co>C��{�ș���_�k��aJ�g�8C��1�*}��i�_�¤�0�]�r��B�	V8ly4(�?8l	C� Z�B�I�^pQ�I#F��ؓ���=/B�	NM*hJ��ϠČkq�إu��b�F{��d	@�������"w.�Q��_��y"�\%N�����m.2�8x�%l�<�y"�یY��uj���$+*M"%�֜�y򧞍�����'�d�E�P��yR�^-�:��@(����!��y�fD:$���o��̣��[p�<QӏU�8�t1�枾P�x8p���<� l8�0�!�D�5�g���Q"OJl[V�D�d�($��]�o�jPѧ"O�\x0�
n�q�4�R�@W�!�"O4�آ��Y ��h"/��
>����"O@Y@�I*���DJX�"O8�P�ȥ~�RLb�.ݩLFt��"O<���.�B����/a/>��!3O���S�O&Z�ƦK�"�xt*Я�>(����':*�� U�=���4[%���&DG�<��O%=�J�*C勺T��)��
HI�<I��.�J-r��7�B�WoP�<��,>h\�,�`���^��g��I�<y�	�89���I�.'}�j�/D"m�ȓ��1'̃' ��Djf 7����'o��4���ġ<A�C�ZA:�0b�7_����7��w�<�D�1��{4g�thz��\w�<�� �]�����I�i�2H"�Rr�<�a�T�&BV�@w��8S�>e��cs�<��N�	Ts\I��.�
�Z8���q�<�6�J:|�9x��މi+�����W�<Q�H�kZ��\+9^$�	�.S�<���4�����Ă [�N4�S �Yv��Z󤞅q�!���(�hʀJ�>�2�S1# Z�!�G#l����^⬁'%�� �l��'c:����c"(5��I�	����'�(ʤm�"J_x� 
}D��'En��*ô)t�A+DӇXAع��'$T(c%#7J��q%FI�L�� ��'"��Ӳ �n���C�w�(�:� �).�B�	J5D�U�۰?(�@�q咴64fB�I+i��X��\�R��dZ��ۼF#hC�@~�;�Y�1���YA�ݑsuFC�e��9%�D�1�z�*��\�{� C�	�)�n����@?F�Xܱ4i�9�B�I�]3�,X�"�
M&�TI
yV@��d,��ڤ�1R�J�m<�!D�Z��B�	�:8�ʆ4q���jج<�8C�	?;4A;u�L�	p���#]�0C�ɮ8�$T��Ñ�)v�XC���
C�ɤ	���B��Y
�x���SK"C�Iz
��$,��k���F���B�I�^f�i��B�'���!���B�8.��ZL�"7�F,��������{�Z��e@�`Qd�ZV��clXe�ȓZ�y��ֲd��y���$)#P�ȓ	p$Q����BJA*�����a���R!i��B��.v��@*�" �C�	�2g�4�3��%iO"�Z�Dθ/��B�	�1�^�Z�F��R����� vB�I&�,[��[�j� ���d�>I��C�I��6`��S�Tٶ�r`�F�u��B�I? ���@~��jPV�#�D4D�<yQ�ϳVw",��@H�F�h�gH1D��X���3.`J��ń�[X�]�6�0D�88�GI��6t�&D���ݻ`�.D�(�3*�7�����A)[YN��D D���sN��a'N�r0H�kt6�GH<D��jg��J��h���P9�|	�d:D��Q4�P�k$�P�N����4$6D��"rKޗ����D�V;6�6��e�2D���Lu�
�����t)&���E-D�@�$��)@���7��&D�`��)D�p�bgF�xش[l
�h�&i���)D� R��QH��Ġ���2E�����(D�� �D���яv�~��E	E�xͦ1�"O"0
�)��c�ԙ:⧋G��Tq�"O\=�V��L�Ă0o�&K���}y���N�\�½C0�ߑb��a�#��	�!�D�*���b�U>z|�t�Ȇ}�!�D�-O���Ei��f��yy F�-a!򄏲6��1$F�)_#��,��<7!�$�	5��QtiMx��h�@�f!�Md�X���/'az��Th({^!�ۃ@��t�rn	�'"rx�'
�2E�F�4/ܥq��q�Ä�o�t��'�y��	������k�@�K�y�n�oh �zc��465!�%�ybN�"d�o� 0
j���g��y⮈+�ޡ[��%*h�	>�y�}�b+^��¸�v"B��y�!�!8p�������EN���y�I� 5¸X��Z�R[�٪D�y���e�ғ����i�m���yb�ζ���� ikK�y��]5X�.\���7c&�倧���y����@4P�
�W�D��v"���yr-�*xغ�i�V�O�uY����y�[�X���qf�50q�Q��y�$΢+����!œ(d�B|�0�E)�y2�U8&�tx�`�	�bV��Bsl
��y�M�&k��y�7i]'Y�v��F9�y�&�1)�
0g�$YrLH��
[3�y��V��ɵg�J
�,��'�yRg��Z��B�$P�/�]�aM��y"a�� �u@�;"��Q�_��y�����=���!����yB��;F	��ಧ�W�8I��yb"�Heژ��cԑx��&���y��,5:��&��+Z��H�cZ��y�Eљ��)�̐����J	�y��T�VhF<H��QG��lB��;�y�숂H�Z�K���7��T[3� ��yb)]�w�~Ի�fɇ;���'Z�y�cSk��	�Z�`��p{B���y���5\@���!�z�[b����y⇂09�rTCA�KT`V���y��F	��|B�AA��n�F���y��%\6"p3���(��U/Q��y���(p]V�@���B2b%`I��y�d�**)�� �  �|�h�a��y"�H�|j���6b�NQ��;�y�(%��H2A�CY���saT��y���Z}Dq8��Q�A�H��@�-�y�$���+E]�	`
�@�g��y2�ǡ�9rqJ��~���󇟮�yB
F�9J�%��b��'�z�т`U��y�*��x�i�Ŕ)�tx(#�Ө�y�Z	
�����5jv�7/�&�yBj0/P�}�bû)[Z�YW ���yBg"�n��VN�)u\"����y�C����Æ�J�i���y2��6)�]A"%Ʋ~ �r�kҜ�y���
�;'� q�x�炽�yr��cn�9�nL�L�����.W�y�%�!#p�Yee#z�Z�@$$���y��'nOX��*	�rh9���y'V5�8\sq�5�h�ʳ��yBaX3H�x��@'"��G���y
� ��gލx�L,��lB3��"O�<z�,�9P��gŀ�6@����"O&�jf��>z� ��&"��P�"O.<��/��$d;���	k�h�) "Oli���v(�#P���W�۱"O�����@�j̘�/��� ���"Oؔ	!��PNI2����	�"O^���h؃r2ai%!PF���"O�ZG���h�I��8���y�kYE�љ���N9��؆��?�y2�R�΍ ���L�V$�u 5�y+�|Ui��!�'6i���5�y2E*;�TU���WU�,��KJ��y���[��j���\�y�Q��,�y�`�'{b�r�a�,q�Y�����yb
^����7n��ؐn��yR��,@�XB�
,[9��5JA�y"���q00�	w�	~�l9$�1�y"�F(1���k{|XB©��yR��0x���SeW}��}2Ć-�y" Ҳ~�D�J TIA�xpQ�F��yr��+}�a��B��G͒)�P�<�y�hCu�D���`Z�DA2�/�yb�ݔ����EKр}��F	�y"���'-�EiCk�t�2V��y2K��l��D�	��8PU���y���"Cqt��3 J� �@���!�y�%αj�<��$$�f(X�#�(��y�O߇E4(�`iM�i�^�P7���y�)1c|�i��[��lੈ��yRG͠��I��[�\�l�)�nU��y��t����;�v�Yԉ��yG���ȓb��k��]\��a��,,�����"��cPC��QEL[+u���I!����2<� �)�M�+z�H�ȓQu � ������\��b(�ȓSA�0b���rj|Pm� ;����ȓY�� ��aʀMPHBw�̜abH��K��IJ��7��'�2�6��RP��)��CӨ,� dNS/���y���� �d	���G�<`��/"�����2n�~�i� B@��%���5�0T-�d�	%EX��ȓ,膙Ӡ�,�^���`ٺL��P��	E�'ɔJFIތm��cab	��2���;��@00�/�-���6a^�Sh�E��!�9���k�p�"P�$�	��r�@ђ�I�M�fQ��1Q�,C�Il<,����K�W�R�	��U�v��B䉞���+��*$��.ҿS� C䉬{�d��������iQ'��B��1�n8*�`W���!�	�B�I�Y3�Q`+�,:Y�L��@Īh��B�	�.�n�;��՞ݼ kTD8�B�/D"�|�6.�Vl�$Kb*^�
`�B�	,]�蓮��UN�� ��ZuI0B䉗S*�T	�-]n̨5-�H�C䉚.���įY��zƀ�5f�C�	�Z�$�@�
ҟ�񙒣����#>��i�1&�%�a��5rP�Q��(R�!�D�>x�eO��[8q����6�!�D1%NqrVj�0=S�-*Ӣ�T�!�dH�3�-2�gS>(B�{l=[�!��S5���)^_d���j��!�� �|z���G�^��r��\��	7�	R�O�R�x���	I�be2_�z������4�'��u(���Xa�����)�Z�ϓ��'Y�?ْ7lŐ 0ܐ�$Ow�x��6D���Ê"e9 �k��N%l.�8`�4D���UМk���
5C1 �p;G�1D��p�@(- ��M-%�&�(�b*D����G�a	~ĢE(�&� ѐ�$D����̲��x���9����!���<��ˋ,k�n�L�F3��a��ɔ��d5�4�D�D6�Ɋ"��,cp�Ť���[���=%�B�Ib��u�̀��1�E��!�XB�I�`ϸYʴlң!*EC,f8B�I�tN����Ð
F&�{���Hj�B�� d>��10dse�1Q��E9�B��%;�Ը�c�O���1D�$��p�?�S���$�!�]���֑Yq�� ��WMazR����Y4�z3�.)���zScۥ.!��sO:�i�C]n����� �,3)!�D�&>�4��MY�^����
"L!� �l~�K�	�"��=H&ህ5�!��o�B�����)�^t�4�O�!��B�q��0J����t�d��Ň�g��,�S�O2��Qb�� N�t����*N�M�AOΥ��&R�t������&�s"O��1�@�U�l��Ҟ}��U�&"Of(uLX�@k��##H��t`)h�"O��ӅЁ-�hЈ�-�]���c"O���m	�t�+�f�;	��;5O��=E��dQ+*�! f�#3d��Ǣ���$-�S�D�'=2T0.),-���	-�x��G�C��0=	�R���pg@��nڈ#3��TiH��y�/¦U̼(�� Ԍ��3��=�yr��[�jm1����@�
J�yRLU�T:ȫ2 S2|5���%%�yR.:-M*��%�_l4�C����y�Bܑ=���aM,u@�'ٟ���3������'��'���A���7-��ؠ�ŔZ�0���'\�b�L!f
���@�7Vc�a9�'p����C%zj
�y�!^M�^�z�'�L�xwJ��S�T�I�lM��)�
�'��`�H/}�,}�����Wr0��	�'�:�1Fm�=^W�<�֮R�Ud��p	�'�>IC����i��F�1��H9����<)O>��+H�T9��A=hwԨ�5��g����	�'�u0��K)F�)�)G�C��3�'e�m`g�0E�L���� &��y�M	�w��i祋�_�Ѣ�@S �y����a I�f��?\�$�D'�y2B]}!(@���#��XD`ާ�y��lUJI�"��}�X�Acm�
ܘ'��'nў��q��T�*� 2iٲa=�eC ��dh<yF˭W2�q�B�C�ț�cj�<��b� t��)a�7a�dx���n�<AEؙz#�i��.0^m�\Q�a�<aB,���܁'��,j�ض�b�< ^CȺ(@��'�ix�g]�'��y2��*A����U�>��@�	��'���'�@�aE�2rw���Ꮒ4#�	�
�'vdq��R�R�_r����1��S�<�Ւ.�-�t��@�>R�g�Q�<Y���6\�H�4�ޖ>� :��D�<i�#�`(0��L���dŞ_ž���K�8�y1��+�L�1J�/�RL��S�? 
����D�?j!��7BDD�����Lx���#�S28A���-9�$Ȱ��8D�|��bï')�����j�d0t!6D�h���X	r��4��|��5D�̚СW��QhC]�n>�ͫg7D��P+�1ZE��"�\4F��g�6D��"��5���"���%��2?q������a�ԫ�7/�͉��ѡg@0
��=�S��y@}���{��W0��qB����y�j�$C����4Kă�-"7����y�)��;��zmǣ
�V�2Gm��yҧǦ<b�`�DB�:��X�w���y](p�(��Q�7f���*��H*�yB��m����1)�j�,A��y��4��!Ɂ,� A�*���O£=�OP�� ���jL�Ю��≮�
�'uL%Gc�B��``���0Wj�9
�'�R)�7-�.)T�٬.�\%C�'��ڢ�C/G���Tn�;(�4�'=�=���V�c�	��.]�-�Ι��'��1ꆆW^O�2��#���S�'Hp�!u�%of���ҀV:<X� �
�'5��J;��١��i�,��'W�"2�ǣxl����]�dcpq�
�'C �;Rd\�{�T9���D�c���
�'���fh	�+�R@��)Y�Y+�DK	�'[�E��h��|AZ�bG��M�К�'�8Ȳ5τbZ|��!E�T}*�'6d�%䛚v�
1q�Jٵ<)�'�X�;�$P!#[8�4 ��7,�;	�'��5i�9y�6��5�1�*L	�'`�ag��{'�U�� T�X	�'�,�c̝�2C�!:�c�1	����'/૧�@`,(u�#�_�~�f,a�'���A5E	w����0I,�ܐ�'�F��B�
D�D�@�D��T���z�'��Dj�L�D�~$s���4Lb�L��'Y ��!�\@�x�S�`s��D�Kю�+#��B4<�$ɏ�mP!�ԣ8�R�k�I�\.@����!��%S��a�ڀRC�@;���w(!�đe�����I$��{WGߙ6C!��;�� L�O48�Y�/�m�!���l���u�Y�=���K�@�;�!�J�F$��'.�� ���0��$2|!�d��9�mH��� ��!A� �rr!�Z;.9r�����:��2�ȼ<�!��Đ3��P
�M�1L.\��dY�e!�@�ƒ4�F��)�����9�!�*�A	&�C�� �<g�!��5*w�,qĀ�!2�6�1�o�?^�!�DՌ=��`�ˆ)�(hx�H�$�!��DB��%yR�	 �J��T��!�$ǣ(~�ѳw�w���o�/�!�ēh�flɓ�Q?46�(�gn޶tC!�D6s�D9�B��A����D'__�!�!(��[�/� �`�[P#6�!��p4����-�*���Aq�Юr�!�d��S��P�B��&B�dU�'C1G!�D�@/lc�AG�kʕ��� �h8!��<^��HW�F>1 ��]�*!�d�4&L}it���Ql-O�2{!�D�*�j�c��!E�FM����<XE!�D@���W©/�84���# D!�� q2�BN$�B��+I)����"O��Kce�4yĂA�6�Ȑ%u"�"O��xu���
{�؃�A�N�$���"O*��CŚ��D��`�zh�t��"O��
���BK��x���hfe�"OA�%M�g��D���ǤY�xM�2"O.(�3��9%�T����3&�4壤"O����E�@	� :�'��7��F"O`U���H���Ð(� r"O�E��	�|��p�R	h�p�5"O�E'gM��ĳ���_LM2�"O����JN�S&%�/�'kP�\�"Ob�Wn[�aj�J$��9,8J%"O��T�ˢ
I�{ul˩3�5�T"O���$ƖӲ�)�*]�
%���u"O�ԙqE=mǸ�8�iT4�T"O�`Q`�pF�, $��8$�"({t"O>Ha$L��(�b�h���NR0p�"O�Q�Pg�{0u3�DTL�P"O�d[ n�+3w�aS�I�lP�"O�� O�'�&��v�3G���"O�9rV�	[���E')��Lu"O�(B��<�<��&�1$�0�"O���E��:r��0��0_y���s"OL7LV�l�0�+"�/gxX�R"OJܘ⡍���j�-�#a,��"Ojq�Ӊ�6| �[b��VfB�
�"O"aJ�Wʍ���W��[!"O& (��k~0���+������t"O��+��	̝�Ɗ��2��t��"O�#Bd������p�扁�"O�[��YƬх@V	t��"OLEY�E\�Rv�Jc H)�6Z$"O>D2���Q[4x�A�W�l!"O�	���$�t�zӮЯO4��u"O��sa��9tjy��-�uw`as"O�mX��KW�����Ra�$��"O��;'ʐ�Y.��� �Q����"O�tZf*� 1�������ce"OR���G��՘Ex�N��~Je"OZ0�B`	-6��os��:u"O>��3�N0\W$	I6��u]���"O"9�&ͼw�����\o���u"OT�P��#op0��3Ɇ�F^�	�%"O05��.��=��*N�&Vе:"O,��@g�d��mwӧ6J�2"O�6��7�2���.T(4p,�"OF	ɳnZ'�B��U���J&=s�"O6Ā��~{�h���,�
E��"O�-�a]�J�iF!-$N��0"ONmK����\��u�WJZ�f>L�q"O*�(�-D�G::|�IN0��6"O�	؀c^ _���Th]:(��8�7"O�-RұF��ͳ\z����M�<�)��K�HX�J4�i)��BF�<�g���J�y�lF�+�Ƞ�KD�<!d�KL|Ќ1��30	�A)�#�}�<y�D�<L���b�ݬ}% �xFşw�<ɶL
�����CK�	b8}X���J�<�С�ml�1KvO*[=\�#��I�<�p��^���!� �#],]C��B�<�1H[)N|��'ة+���q��x�<1�!Aq�I�G"آ*x���Mx�<�栃<M&.�����s����Yr�<� DhS�-/�l�5�����"O X1M8,2e��f͒�~�r�"O&�XG�Z�j��ؒhN�1���+"O^�ɲ���a�8A!��pxL�R"O��&����h��ܺ/O� �"O���� @#;��!��F19 ��"O�̈ ���L�
��@E�&Btl�W"O���B�F�`4꬀V�M�y:4�"O��)��B�����$�>4�M�"O@}�I�P���i��εGO���g"OM���4E��!y E�EY���w"O:��%��7Z��ש\�MgA��"O8L*� *	��ѷ��_^	"B"O(���(U�ߜ��1"� ,��"O>��ΰ.��ᚺ*3\9%"Oz@�Ɓ�/\�����A
b���"O���''S�e�2T !+��=O�=#�"O�h��@�B"b��ţzQ�TR"O\U���r�JxP��Ȇj�2""O�������.\��	֘H&n�c�"O��BcCH�D����
��4�"O��)%$T04٨�c�� c�4�8q"O�=�rdRW�$-y5ƅ�'vx�"O���U��1iJL��k�;u�9�"O��9�� .�&�h�Sdc��k�"O<`+f����<�@�/JytH��"OX,酃��F�
8 0)	��  7"O,l"�Ύ$%(��B�֐j�"O�D�,�	��Q��C�m�~dKs"ON���I[G��82d��HI;�"O���n 7u�D Dӂ��`�"Oе5@�����/�/~�i��"O�#!ێ[�����V�@I "On��LϽY?p��D�@2a���`�"O�DA����:�4����v�y�"O�{���Y�@5-� ڈ��"O��2`=�>9yt��{ֶL��"O�]�7T|�3-�$�lQ�S"O��j��E	-�&=3�l@X��"Ol�z�n�0H2��@�01�I��"O�ؠ0��j�JLx5�J�S��l��"OZ�qD�>�$X�/��;��a�"O�]Q'A�� �PU��\�-�|��"OH͛1�H7\"!���QW�|�x�"OTP��Wb=��3��SQf�#�"O�XC`�׆f�
�*P
B;��BE"O����\��r�1C#�؂�"O�ś�fL`H��Ƙ�NAT�+3"O���7(�D�ufܙ%x��r"O���WK��eM
� P�̩8/6�a%"O��K򊚧U�*AjO�?�D�A"OΝH�A��߆xJ���B8\�"O.��0AG���0"*����5��"O�ͺAD؀!1�(ҳ9��F"O����$�R�C�'�2 8�y�"O��R�P$B�t{�-݀�1��"O��C��nJ�P# 
�*��zP"O2SbQk�@eC�@"}�TP	"OX�HF�4;��`vc����J`*O���N�,:����nϰ_���
�'ê��qA[� �l�ڰ��*Hc
�'�:�Yt��v�D�ǫi0!J
�'FtP!蟏m5�G�f�$MR�'؜�H6k�V��<�1P^ ����� �]`��C��`��*�;n4��1"O��c�8	�<�ACR�i\�#"O��� (��|��A:1�t�s�"O�)���E6'�L)c�
Y����T"O��5G�(Ђ�:"C+NJL��U"OT,:� �	{�b�A�D�%.��"O�����&�,�f��{h� "OXy@�g
�

]��/�p�x��"O��P�g^�%ƪL�`U/j�n��"O���`��Hw0�2A�ҼR���Q"Oځ��j[1(��蛅͓a{��)�"O�����RG�6���R�]p��*�"O�a�*?��!Q��Rp�EzD"Ot��fٌy���ZYW��Seȕj�<�q�&2�j�җ�Z&H�"���oDM�<9�� h`59f�]��hT��e�I�<��8I������L�������OZ�<��Fr�y�h&�8��r�
W�<�
E(MR��ք�m�t����Y�<��T�	N�@cu-��b1.)�r��Z�<I�+O�J�^���Nԉqc�=O�X�<�A.�iX��`/U�w�[V�<�lӛ'{ �keh��30ɐ���W�<�с��]O4X��Ĭ}�v�8c�CR�<���*p%�3h2YT�ypR�\D�<q�)]���Ro��-Cd|�_�!�؉3պ1�Bk�%����H\�]�!�dƨl&��F�Nh�]��
��!���T��Qʄ�W�c���S�F�!򤂫8���〦�:{6�%dZ�a�!�dG�:��}"#�_]Z4���K"B�!�DW!��QK�蘩2�,"���!�*�eZ"�ЬS�%P5/F� �!��;{�>�S�$R 	fF�<���"Ox�Bc�˭DT:�����`�*���"OnE�eN�>������T����0�"O|�!�kF�Fe�݁4.زTH����"O�M	�kN�h�9җ�1E2�"O�ГvE�3[��G��ED���"OZ��� L�{ޖ�B%�-O
^��"O*hCd�H�>3�tU�� �@ ڳ"O����
V�Z�4L"��*f��Y�"O%�rg;PLak��_3P���(�"O2]����Q�.��S�L-H���w"O0z���o�Y2 `��'��H�"O�Yh���p�`��űh�$=�"O23�T�G���� �v��@�"Ol5
�Õ�Ha�nA��}�W"O��RC��c%
�B�L�w��`�T"O\= V��m9N�� �Nl�{@"O�B�� �*.e:��%���"O,Q��� #��(cGBЁw���R�"Op�`�f�
Vhz`+Baۤ���"O�`Hè���L	��"�<	Ɉm��"O�P G�@������G��u{"O�Sr��a3�|�u@�0h�|�"O���˲`��� PM � �s"O��@��J��Vd�t��sg��Z�"O2��1`,<�j���I�TTM���' �͆�	1�<���퐑zl�sS���"�,��d#�DC�N�
��끗O�8��D�!�d�&��PI_��y���E*ў$��llN �p+ �?��C���RB�	!V���*ؘ�2�hV&Ur�C�)� �T�T��S��@B� �c�@I��"O\m�c$ �#HL�a@E9$l:��V�>��p�<u(v#�L�0i%�%�v]���3��	�&RJ]�� ��^@p�mKGnTB�	�Vi%k�G<y80��F�x}"?Y�h9ڧCr��n]��=x�Fχby0`�ȓ/#��чVI�>}�Վ�P"x!�'ў�|�rA�(�xE@C"�"Hʔa⥃j�<1�#{�f%�&�*5eԝ�`�e�<Ɇ!�W�Z�V �"`Vt�⡑j�<���-����o�%,]Zy���a�<Y�[���(P�)�$8-���V�<	Ć�9V䡊p+�b��e�l�<9��0;�d��D�,8��T�f.e�<7E�'"|qxfES&>܂2_�<yDNc�T��D�UA�\���R�<��EM98>h�ڷ�� .%�U`�(�K�<q�FO�!���R2���etd�ԀEF�<10�%KAf��֋X� �2�fIW�<����2�&��F
 �ݺ��Q�䙸�0>9�E�:y����@�]�Ђ�@�O�<���G1_�| ����_����ia�<a�#Z�Cw]y�D����*�[�<�р��1D4b��1���2�^`�<a�,MU�$�$�� ZhS@^y��S�n��OQ>��"nT�8��!��F~��h�A D�8��@C�	����pπ���B�?D��Ԭ������@
[ B��<D��2A [B~���$̶xz�xG�9D�(3� �l���Ix@�GC*D�(�%Xb�dm(����馊)D��Չ	�X=\y�g�;K�6�Pԅ-�d+�S�P�tEC��8RsB-4J�7���jϖ��d�[�<$`��tA@��>�דa�P��vB��HVM@C�	?L�❇�5~Ͱ�h�Af)�O��V9�P�ȓw:XL�p��
�0Ơ��)�B �ȓ6K�t�x�ʱc��>�N�iƩ4D� Q�^�@8�dCg%ߨh�U���3D�#6H�7)K�+��JM�@1�&1D�t2�_'5��ꥈO����q�.D���n��,����p�N�z��5�2D�d�ʋ	cs��q�W������1D�PX3���5�ib��ְ�r�� .D���L�9kW.)���U�6t��Q�*D���U�O�I��(��R	N�X�(CJ(D����O�4
tJ�M��w!�m�s"*D�`XtBSG���l�q�f-�%D�D�1�ݘ@�F�2��K"�l��1h#D���$-^�1�f|r�N�5N�T� D�TR�`�5�9����'&/�@`b9D�(�!��s4���D�2cH(<�d7D�@r�0y' %C3��(c� �@$m5OHP޴G�%�<��'A�j�t�aUkM:W�&�aTK1D�,+!��*sրtZ3��?AĔ�� 5D����J IF~�4��T�����i4D�����W;x�tIڱ4ւ�"�3��0<!dB�n��M!��.o��� �F�m�<i�n������#HW�=��2�,�l�<�!�L?I�v���i� ��ܺ'��e�<�`�?S��i��Y�8���ⵉ^�<�)�d��\;RkV�Y�ػĢq�<��^�L�������vvų$��s�<IH]&5�	XR�9R�V��pJ�s�<� ��h]�4ܴ��w�L�6��"O���s��$M<��'㕇7�u�"Ot������ ��@Ig�I�"O�db��E�Z�B�w����y�"ON"�hW&?� �@�nJ^߲�S'"OF!kB@�\��Aa�*Ͱ��"O�Q�K�'L��(rW��;k��]�f"OH�#0��#�89!�F�=���c�"O��� ��5Mq�LՎZx:�¶"O�T�$�>K `@�F�|Y@��"O���G! �TD1Z�F�����5"O�����N"N i�<�,$�"OrW�
Ҫ�j���Hd���rU�<!��<rIds6�Hl�����Ih�<�ˊ�>V��bnz�z�`sCNJ�<	5)ˆ8nj�����:Ƈ@�<���	�>�cR��*8P*]ڀi�z�<SC��	����M�j�T����_�<y��͵R�.8rӀD	sq��
�˞t�<A6.�"K躑8c�K)aɦ�B&�Wr�<Q��7���cd_՚H��"�k�<��!ܜv�a��܊27�Lҡ��c�<�&	Ҍg����˕�"��TQ�^�<y7�40�Th	Ӵh<�ӦE	X�<q!	��{�eӣ�c��L;�dQI�<����)��܋rNE�
��Ӱ��B�<�S,�'Ft�M�e�A����B�<��,�0}쀀+����}�,䋷��F�<A B�_���q�	fI����	x�<�J�[�M{bn@0S��y�$L�<��(��o��kL$x ٣"�L�<���$r�v�`�ɡ*�t��T��^�<��#����IQ�̞
������E�<����E � �& B�gc�T*a@�<��4gxX5���FE8��fm�~�<透��y���s#ڢ.�V��h�y�<��R� 8$�`-	;Ğx�vfN�<a�B�`|ȘT�3�� � s�<�$l	�G.,���\;cL����V�<	���S��uK�40�!k�#�Q�<)���22����@Ѱ,�)s#�YH�<I��G �x���)5X�rE�E�<��@��^�IyB�ɢ6"��;��H�<ɀ �}�I�QH0����G�<I� d�^�� �S
�2�JS��k�<�Gaڑ?�<������[.�:f�j�<I��!�(5¢Μ/�����c�<�Ǔ%m/&c���<̞�z�I�<��`�bT<���ޠ��8E��y�<	�!X&{m��f�|NP
2�l�<91 .O�$mS���'2ڮ��K�g�<�"��N�6\�5ծ!"R3�@{�<�3@P�&P�A��"��	#l�s�<��,��H]���(_�����n�<���s�H�� ��1��(���c�<Q���2>�JE�&J�K��q(�e�y�<�R���`�V�*�Q>�V�г��M�<q5c�#+%H)�A���`XP�����F�<9��
X���-���#�m�A�<y6!ُ`Pf9�W-{")�w.^r�<AVLC"T��$���0A��P���Vo�<�f"��(���֫">���l�<9�lV9m���#�I��t�;V�S�<���K���;ӡ۴ ����3�L�<� N��(E�J��Am���}��"O�9���E� ��XY�+�18��92�"O���X�w�|1p��A��!"O8��##]�y���c��$wR�S"O��k�.f"����$����"Oּ�w�\5�NL��֍}�
��$"O<�8�L9t�����6� �"O,��v�
�f,N���E�2k���)�"O~a�i֝0j���r�S�x��"O�ɹB��U4�`r�aAK�p�3"O�-�7���h���JU�[�2Ӕ"O�4C�@����"#E�x�V"O��[eȅq�HU�!�Ӈ6���jC"O�Ix��M#:�r���̤yM$#"O�Q���Pq
���r�W#(��h�"O�H�G��y*�#�O"J���Ҁ"O����xwb|�Ak	�$�PU"O-���A8���K MԐ�1 r"O4dŎt&��P�	*hz&!��"O��0�"-4��T17�K�1l���"O���R`�1�B%:�.̿*k�P"O�|�\G�i0�nƪZ@ѩ�"O��:!N���iIw��- D���'D����瘸e��Q�'�+=�pb��$lO��4���ʊ/�Na�cCڧ�<��=?���ᓥ�nyT&[�/�R�Ώ=:ΓO�73�S�'(�=��
�_I��jO��f4���$h��ɪ_ H�1/AZK���>�2�'���� 	F8As�B"�:EZ	�'z��C�9˺`#Ю]^�p #�#D� ↪��GR��p@��6(��z��,O�#=)f(�R����؊!�ʥ��@�<�rb�	�F��͟ [���`�%�{�'T�x	�m�FD�Q�8�.��P�:�HO�����IJ��Q �T�dc(�bv`<>集�'��O�Q¦,�	,޴�!��<�ޱ��i����޾t<<��f��_ �'DT�m6qO�=%?�PƁT����5<aIӶ�8D������wl�Q�gAX7> e��#1D�PJ��\�p�@�i�!S-,�ވ)ba3D�$�2dɥ �����D��o��tz���Op��0>�Gĺﻒ���ZƎ�A�����I�<1��OOA������)\�))���H�<��܂o�)p ιD!�SG}�)�'n���`�u�4���Z�4�\؄ȓ0�����¾09z�`2�\61S�9l�B}B&\�<q�'xQ�p��_]���:������=�Oj��)ZPp ׁ�)@�p��YC��	�o#Xl��I�B�RY8�L:���+���O�?�O<9K?1ʶė,��+6�;]U�e3pf8D��We\�8�����OOd	�T/1\���<�O�6����7n=�wn_N�>��'����-��8嘕�һD����޴�hO?7M�0N����@9�$G� ���d+�S��M�"�ʹM���"c-;/�貒�U^�<�U
N�RTx�6J�|�V�ʗG�q?1ش��>a'n�?3
$���@� E�Ng��m�g~�a_�u�,����G��VIˣ�yr��&vB���D� ��JS�[�yr��*e#�$��N�鑁䍭�yr��+YXX�çd�6H��� #�yr`P*V뾑�7b�'�ĈV���HO���ĕ<8n���v�6�l��,ե	!򄙂LI4��$�T�J�R�;ū�1E�!�� R�Z�gӌ�,�0���)���!�'�qO��PDn�E��U��]?�|��"OBp�u$�7�d3�*C|�>�Q�"Oƍb�-_9RRKs�Q�t���"Oȕ��\��Ha�J^-~�����$|Ӕ����:�	���� �䔚AMܺ[!�E�8
��c��U�e|ࡊa�ۛE>!�$�?+|�`⣆�td�B����K9!��_>��;tm�(JO��xV�φ�!�$'a��q�U��7iAD�b�j��a�$0�D8?%?�'�Lk�I��@A!�˅in:E��'���B�#A������?k��	�'��D{a���K��ꡣI(D\tX��'h����`*��x @F7uI�����R1 HB�I�r�jAz�ڌ&�dâ�1�B�0p:F�H:O��ԅ�=��C�� �� p'%G�jo���%�H~.<B�I[�5����%-pxB�L�D�nB�	�M�zT�Tn�]�D$8u�M�N��B�	X���Ȃ�1,\1�Jq��O��=�}ڄ��<��� A�Tbt}�Q,L�<!�����Jp�XO�R0K�	�|�<�Tb\�Ik�Z� ��G�P��&x��Gxb/�%�>Hj5h�y��Is���s��B≴=M$'&�1�¿ۤC䉭-ڔ`�B�ńk8�1+�A��`��r됽#��o���Gj�� ���Ey��|""m�m��,�狂��Rm@���V�<aE�ζIs��7�&t�9(F�I9V��O ��<���ن`F�@!���q�rO�<	U.��g�j0���z��[WI��P��I_���O�fb�R�n=y7� hd�5��']��3�����Tr'*xc�A��"O�`���E�I`�ĤK��XZ�"OT�j����$*ǃT�.��,(W"OڤKc�6"N9�����T��V"O�%��Y
�2@ �'S�@�LH3"O@=3,N�>�q��)Z���0���F{��	D�BXz��㉐t���:�2(!�d�*#hB�@���c{Xݡ��Ԭ3�!��8mⴠӨ0F��)�i�6�1O���O%^����@*�,N�lHI'C�r_!���(��D� ���t�(��S�Ñb�!�d�%C���v�����@Q�{�!�$�8Z[f�>G(�!0�'E�!��P'!��U���L����Č9�!�dۋ?���R�U,z�N���3�!�JJeBIi�䁿C�d}#�P�y"�I��v �6"#!�J��jP#
uDB�ɜn�D��	�(hl����B�1���9�m���f��'��!$rlB�	;4 �#FX�aD0*"�B(�J�O\�=�}���ٸ?�l@(�L��R��x7��p��4�S�'7��c6C Ϻy��'s���?A	�}���G�A~���B�H�ȓ �j�A7�_�z!H[�����ĆƓ襳�d�
O�tX��nCX�^���'[Z<�3-ȉ	A�<���ӈ}�P�y���'��e����=��`���8r>�(2�y��)�S#r0�zu�Ü^��%�F~-���)�-��"kIP�#���!6���Fx��'&��2C�.7S
�q�C�8�|�(O6�#�S�O� ��)^�c�,�?��,����jh�r�g'�ő� � 4`���S�? �%{PDX.�q`�<jX�q(G�$G��(O�wn6d{��Ék����#��x���|D{��T"�(_31"��Y�64  ��'9�HOOfc�`S�O�k����ʀ6GR��o=D�<�%((GV&�� o]��*+7�~��C�ɬ9����u��`�|1�.-�C�	1
�r�#�:Mar�-E�Ȍ-�!�dA�N8r�B��,�X��hňI�!�ă�x�R!B��� f����ЍV 	�!�d��),�/N(��I5lW�+���hO�Sy�D߰%��]���ٷ)���ۊ�y��^�^5������!��L�M+
�'��Au�1FT��)��:�z�b�"O"��GڏVwޡ����x<u#�d�>a���հ9DlyeŎ�
�t� ",�V7!�$K�w���pe����̘�ző�4��	$p�ɇ�I�#�����Wk_HB�I,\�H�h��?h���zU�ӻ��C䉊�����A�%N�ɥJ�3EG�C��*8��%y�mZ*Wc�<#�IM?kPݛ�'	5�ɓ���d��ʗ�6�y��'�NQ`bX�H��`�5(	7 B�Yk����dA�I҄�P1��0�8_�(��g���&$KZ�ؑ���J>����B�>hB�'�J+ �,\��n �&Zn��ȓE)|pr�ĝ�W�`QI�'�*onńȓ-�X�RNU�7H�r��ܥ8ΐt�ȓ�r	âf��
��$ �F�ȓ_BY��EMy��!���ŹJcq�ȓlH�ۖ�\���jU� �Lą�Hm6�@�B~��Ta���;l���ȓ ZV�ʳb�Ȟu"`	�A�a��'��xW��}[pIr�Ƃ�O�ۅ�b��e�#-�{��q9�a͊S��l�ȓWj�a$ˊw�@ a#i(Y ��G=6y����c�l���
ROu$���hv�" @�iuj�8��RM����y����̗"b���DiO�j�0��&�s� �2
J�R�G%�vp��/@�;�(Q'��l��V�.��Q��?ޘɵ�S�i2���,��?|Ʉ�3q����V a���g�?A� ��Ϟ�p�K�\r�
A��7,*���t���D�Q��mv�ݵ����ȓ
��Q��D2X\ʤnF�2���G��Y��!�
�b$�@v&�ȓ	����`'ŸJ��`���[�������x�R]�QÌx��H�W<��ȓU�м b��M��)�-�5}�`�ȓ���æ��7k��ɲ����FU4�ʓÞ\"�ɘ�1������l��B䉚v�A��]�y�P�t�˅lbC�	D 2���R"���ѓ�
E(�C�	7!�,TqQ,T�2�hr���&@tC�	�@5(�)Dd��+r�M0��O�O�TC�	�.���hF/<"~z]y�$�%(C�I'U���X�b�-W�,@!mșnD�B�%Vr�*�.�
(*�(�  BnbB�	��Rhb��@/?L#c;KFB䉆|��0z����q<(�2C� [P�>�w�� �0b!B�.<�x@�Dş�q���"'���q��4�X���>D��� f��b�lk3�(/��aґ�<D�$�F�M+�LQ��$ 6V���K78D�� �mµ�����(k��	�7N,D�� QsV��1!䀈�� ъb%��aF"OR�����#D��5���7(�("S"OhH��JV�������8L�bĺ�"O�h��M;Z���Ab͆��z)�"OD�*���=)����O�<�zy("O�D�L�=}m����
Q��t<�"O����	U�tSV�A�M�@�@A"O��f!�.:x(��H�=2�f�b"O|�X�M�7a*Ҭ���W�}�J	��"O��÷IU�i �����t�fQ�D"Ov�Z��|�BP���W�6�l˒"O`h��dC/Hf.�4F�L��8��"OFl�f ����}8@bJy�� �"O�st*�L�N0�K۩\P��S"O� ���6�cu��rHU�c"O� ��Ǌ3u8H�
�E��)�"O4����F�R��3h9*�A�s"O���E��[�����Q|��d�"O6)�p%E��4h���	E�੷"O�Ђm,?�XµH��f���"O~]�Nї4��9Aߴ^�(,AU��Ӆ'�n��)���M(�X~?TW���!��:+���[+�d�$e�Ӈ�1����,�	��H���3t� ���_�d��Q�d�%<B�I�G&�dڢ�D�@n�Yb�K�`6���IP`��
�\X���׳p&yGKWD���ɥ,�v�2�X��fZ�F~r}�-� )N�I�=D�� ���Ux`����� |���'����|��q��KTӫ
�:P*�O �zZB䉆{D��uJ��=��h�o�	,t0��Hܓ�>�\�,�`�gIiy:��	�3����
�>��Ăɢ������/���	-O(�$��	�7>���埒m��y��L8�B�I
V�#�M٘S]���Ɵ|��B䉥y\hW)�_�B����M@�C�I'b�L����7Z 2�AM'9`�B䉋�6�ا蝰AD,�(�j���U���Y@,X�#-�qZS��-=!�D��Y	�4:�Kft�YC���.2!���X���A*�U�y��,�!!�dѽT^^qzg��9���RK6!�$�p��ɨ�'�1gsF����+X/!�d�6"�(����M?&|.��K	�!!���j��r� W�L��Ѫ�t*!�$�p~�[6��f����	ýj!�DR�8dЀA&��%6�ڀ�)�X�!���xb���;3d!*�(�s	!�Č�D��,�E�U�5+�䛡�6�!��P*.��k��Mb��8珑�l	�'c��0��1�)��Y����'K��x�`�/H��C�I1��s��%<�@�7��pژ{`�x".��<�9�}&���B䈢U���GfC#/�xh�3G0�O��r�HT�������8V^�3�#D�&&�a�/8NY����I����PD�Є/c �:��ߊDZ�"?���F"X�,h1S	� g�R �O���/�9$���U>g+@��'��p�c�!>�:CB��7�8�i�'���HW|P�Q�Ɍ�|V:�~��nߘ+�*�"���#O�Xt��x�<ٴ�D��v|�6��$uAz�0B%�Nm@ �Kg��q���ȮA��K?��b��B�@Y�Xヮ�`�,�-*�Od��Fe�2nN(JV+�|�y	t%^�T�b9�6�� `�­��A^�AV�{ҫ�K��k�C�F��R�,pm���@z�" ��L$����ْv�ı�'R�z吢���I��QRq��!����I/Z�Z���TG��̤8�vtӶZ�]����Qb�M�"+��o=������.�T�%9��>�2�J�,\���������R���O���3m]���)P	�g�? ||k�@%V��ڭI��L�e�F�T�*�d�Z{���dω]*����'#&�P��F}Dl�ǂ�#pA�ٙ���	��#E�H���i�X��k���^�C�A<�̤Z�.^" ����`J�;S�
,�C+T����ݨufH��3o0����=j�����ǂr�¤!K>�a��q�ЌA#�Bk�����O�Q�dʋ��n��%�W�[(�PRw�R-��d��s�T$�L<�AbX�v�`	=?� �&��m2�[-�|H�L���lRP�Z� ����j��:ô��P@��H�4}i��Z7��0��B3;�}���:}%b~��4��u��$gr��D#�<��n�#�B�pឤ,Y�e�r�A�:�f��NT6�Q��ݴ(����.�(�u��D:�j�7@��
:H���%Dj��*�M��6�J�� a���`�b�y�,�c��# �$��y刞R)H,�Q�ػg�"2j�U���'Λv(	�BrF)�Ǖ�t��S��u��Aωv�dL���n&1O��Ξ��`aa־C#��@A=�BD�ԅ�<O֜��c�Q5^.�Ђ3Oz��T͉��P7]+��'��5	E��c�ӧX8b#ז*<�����Ž|�����@�NO$(��K��S���IN��g�H�X4j7
}�9�a`��![rQ1 O�c����/K������K�w]�\����>�܎6����S�W3t�Yj��"���x��'�<)cu�G�'�Dy`R�]5��'ML��pd�f*�Xa`N"k�,���A^�0�䨡�C	�|��!T�;�*j���y�U�xԘ��ٹS�� ���U��r�T�Q���5��I��*C�S�]�ƌ+cW��4 A'	��Oty
�L�AGZj�$�f��1�><��i_�������<	-�o��aZ�����	��$����|�iN7�R��]�e����o��� M�7�_6����h4X�Ӏ�56�����B�I����d,N3]p�Y$�ā$��_t�]���Zg���Qi�>��䙗%R�W0�<a���Y`̸�A�>!��A+�ʈ��"�I��1��);�̼����*-/ C�I�4X|��ڳQ�Z�X��� "�X�B��oˢ5M>E��b
�9Z�}:��1'���rP��y������.MJ���L�8���'4�}yr"�n��Z[Bl��{Zw�(]X7�!��k��U�`f:�J�'Y�%z�KM+e�z�e`։Pb�A!�'k^9�Ð,�ɧh��l�tFZQx�17�G����F"O�x#,ʑ BT��P-N�V�XA����tƑ Y�8�`��'���7�ܖ1��)c���:��\��r|���PM�=BdV�2���4@�%�B��n!��&5�̈6kO'�Bѣ4fD�!t���/��h��!Dܪy���>a�A�N��!�b�$E�tH���-D��Y$&شR�<�(�C8���ZQ#|�DՍ�	6@����>E�$a �UG`4�E�_�s���)��߿�y"/;i󢍒Uj.noN4��^0��䔝_�Ƭf혼�p<���%W<|a8�*̍>pD�p�l^d��0BV/�rG>��i�
g���K��Vp��fБZ���Ȃc����M%k���sD �HW�I ��خ��t��պ�,\h��'m�>TH2=�!�䇇����e]e�	Xw�׀5N�d�-� <k7h ��/z�d�T/E�E�UBV�J�#+nB��.x���W��T2�mP�O�{<�\x�'�T��#?���0b�'Z�-����F�~9r3,�%��T����¾]~����-��v��Lbt	�2a�b�j�1(�C�I�l+fl�=}VQ�N[�B�cQ�	��j�92v8ҧH��Xɠ�ֲ�j4I`�]�_A�h�'"O��w`J2�6u�SIx1��	�	*}�'��"�vĩsd3����&^�1QT�_2.�Ɂ�Ф �a2$�.H6��2��cXJ�9w+D�3��i��
-f��H��I�o��L��D�)~Ex�kI7S��"?AǇ� ��e�h"��G� ��a���C�Ӥ}`�Κ,xn!�ԭzP�E�U�~���Q;F�I *֜�5�Ue��S�OLp�"�$`�t�{�͖j1�Yx�'%$(�PF3=�^���N^�2I���t�>	A��o�۳���}"G� \�"6k���	(b�ˈ��O�`r4�˃��q�pZd �/7a���K�-U�ʐ 1B���Z3f;�ON�J�NӷE]�Ժ7�Z9L<�H��'�0ms��N�z��{�n��]4Ӏɔ*qiyD�³�!��2#FIr�'T�SbX( ��<���+?�J�:���|x�OH�Uf��?�O�䋁�]��0c��.���/@}�AI��5��H��L��(�F��X⊝��HL��HO?�$��A�Ld��*$�\�y 
�qc���3��#L*�@x5�� eaE`KJ~���������O�����/8���v͚�kH�#�I�;\6M�ܶe���I���)��f���O��#���_��[�h��T!�dx�2}Y�'�M�>ıfl����I"=�:XZ7aO�a�8�Gz*��q`���eg\)b4oJ(���h@�'R&E�q�W =�;�J�X���#�ߘ} �X��R���"~�Ʌ�KƦq{Xm��+�~p�9B�k2�Į��<���
�C 4�zX�������#�O�pzJ���.OL��m[<}/i��N-��'ڲ���"б!�ɧ����ś8!�*a��όY@p�hH�C��32�2�89ׄZ�i��9Z�N�5S
=��<?y��j��&�0T[V�#tB�ӧu���
"�%#�˹���3���y�aۉ����CE<��yQeV����"N�y��+��)�'�%H��Yz�j ��	���^��(q�Qc�h� �tX�1ĒJ�F$�J���d#�&��`L|�>As�A�3�dD�K��P4	�d�q؟t
�� O���"%�Ƙ.��[Q�0\�����I�P����X�:���Y��ņGoƄED��$�0rK��cNO�����-���z{����T�sԐ%O@�s�|B���T�y�i�fb�/�j���C�VhV�٠�O�@�wN���P�J�"}����[�fl���KX������[J�'�za{1I�2�D��KJ (ts� [�4�1s��!��,��qzZ*A���'��԰�i��E4:8؅��.(�2��_� $#C������1+�5;Xl�`3xrPs���)X]�H�Ov|[�A
�0S�e�*?���c:OP� �2sRXջJ�<�A�e�qOJX�c��h�Q("����AY�'����˱E"&鱄+��9��"]����f��y�ꍚ/��t�@�I������C1�O�i�e�3P`��Ԅ2��,#��W:=s�h��3!�!�ݐ@��y ^�2u����䃝NP�9���z��:K�"~�C�6�qwbϷN_l�!bN@�T����<u�Mk�h�'�d���%]֩�&�|@��8����*���w-�;9�������N�|�l+2	���i�ze��(ιt�IqCM�!�$��'0✊�oY6PC E�Ca=
k�q�����-sJM�����m�5���Q�r��5�X�0�!�D����L�v��!T��2���o�!�$� j�}C�b�"/��ҁ@��!��A(`�(ij�e�+?�8�������!�$G3$u��9æF�q�`�����M�!�D�7#R"��R�yZ���!�$ !B�� zn�9��ӄ��8 �!��[�|`|stb��tφ1���؞Cn!��$~��xQ#�;|��L�+�@F!�W�AZ�-ڌ�x�QJ��9L!�Ę�?���j3���6�Z6h��.�!�JiO@aH�&f������S�!�$�5�TYXB,�{Pjњ`�G.�!�d@7+�,P�7ꚬ 0�
�'�!���&b�I锧�8c*p�8U��!�$�=)pB�3����4pTQ�Ɣ�|�!�
�X[E���
]��u��e�!��@}t�D�O)x�*��P�H�I���dTj��xBi�"928��d�yҌ�,srVݡ@N��;=H#-̗�y�NO�|��ai��K#db���y�Qtv�e��]��8��a��yF�I�25�c�:q�X�k�
�y�Dݒu�L4�v	G �t����љ�y��E�>xt� ^.�'�۞�yR!��w��X2�� �3�"�y�h_-6��yr���3�P� �%��y��Fq|�v/�
/��!	�h��y��2	�1aĀS�7)֨��S�y
� ����c�_��=�@FR)5*d�`"O.xCU�I�d�h��C�=7�<�"O^�⌙)7��H�sB��(H�T"O�@�SZ�Fچ��f�q_�h��"O\Ċ�i�'�r�v�Y�q_T�@`"Oz�@B�9v��d��E��z�����"Oh	��ND�2>��
��d���"O�D�&�%2r �f�бF�6���"O���R���q�H1��K�uu��*r"O$�c�h�<��j"�ͅhl�y��"O�@ӱ"�:SL�CG�1t$9�"Oak`�2>���E�p�^�7"OR�
��^0^E
�R��5B/��s"OhxГA�X�6Kۖ&�K#"O$ɣg8>`(�qC�Ǩ<Ԙ��B"Oؑ���D4b����ҧ�+���2"O"�kuK�^��%�[�4��@��yB�_|���0�	�y�h9�����y�<P�P%���r�H�nؓ�yO_ |�<�V�i<�dit���y�+���͑G��.pD���Ɨ�y�~
�3���o�ؐ2v�y�JݑR h����E ���
�#���y�I�_y�¥��lxS��]��y%\[� �6�36��p��M �y��N{�*����%,uڭk b¸�y�� u@\d��NN/&����Ǚ	�y�F͝����!B�E�E����y�#�N�v�;W$�1�L�k�����yR/ �6����Ҷ!��K !Ρ�y��,z��	D�=�0�����y�A�Q�V�UD��&Q��#��yR'V2I����C�Z1�A����ybm��Jy��I�|��_��y�"�f[���]�rOx9�����yr+�&lW.�z �T�ZuNp�����yb ޷jX�1��Էbl�@i�y,HRd�
�@�b=�EZ�cG0�y�GK�X��9�@Jϗ�� ��mW��y��A{M8�v�ȱf Qq�H�:�y� Q�K`8�"��:S��Iy���y�������R�\=G`,�b�	+�y��p�@��/�m�-R�T��y��I�5�0Y;V���ap`h�5�	�y�ᘉj&��pA_\h5+��T��y�hŏL�:���+JP?
�۵��.�y�p��1����M�e�t�� �y�(,ve
Dx�(��i�� f��yR��)I�=zW���Y��R��ʮ�y"�S=T ��r%Nٳdh��R�T�yR儠^��p#c�'\��lQ����y�ƌ[�D���HS�f[:�
$�B�yRH�%��@�� ��X����y!Վt4�#�"�r̶�@�*]�y"d�ɢ%�MO�u���W����yĒ-e)��â��.�<�p�`I4�y��Uc�	@ ϑ�>��07 ��yB.�=-�v-c�bڱ@n"-�Fo 9�y�	ҿY�"QAQ�$I���H����y���]#o��l�[U��y���_1
�yq�E�&͊���AJ��y�~�~��c,�
n4`���"�y"��A�� ��E�u���u!���y�bN�U5�Ma!M2`yİh Fа��x�� ���c>"�~@1�k�m�:-z� �,P9���	7o�0���.(B4�F(�K����:.U�|�'�0}RĜ�3p�:a� C�N����Y��y�gM����x2E6F��x`��Q��� m�z�ɰ�M�=�a��-m� �w�\'v
 ,�w���y����P��� �N��w���I%9�&�M�8&:Oxq��')�@���*dJL-2�!u�=c�'|<�@�C�P���B-�qقj�	x``4��J��DI�$W�@%̝!��1gP��a,?1c �'c�O���H�>�Q�Oh���C����G'�U`8�X�"O�%`v!�V��t��iE`l8�j�>�0iӈ��L¥�7��S���d���w��*s��cs� �vN0qԸ\e�9ғ�b�)pg'���1 ��P+�>E�ոp+R���Xx0�E�b��'$�P W-�j�F|r��1�
���D^�x։JB�8^:�9�P	{N�O86�Q#���;T� �Ɍ�V=D ��W��IT�D�&B�P����N�r����)�
���S��P�#�U)|���_ {�e`���;�X�'�T�P��[���$��@87����d.}���d�&p�t��s��xp�|�A+�� ]�ɩ5��[�$���+}r�H
�q:��.�閑v)�dR�\@�N�/6�-  i��Q`�Ȼ3;�xr(H�@h 0[h��"t� h��m��Z�GS:_����DI�V�.��V�����?isl�)O[yP��Q?z��T���7�h��D%�fYӧuk�)�( ��(�}���NѢ磞k��%c��S�CxE��"O�ió�֯7�"���ڢS���B<OjV�r��U(}��4�:�pK����ӥl�j�<�Dy$-C4P����"j�H��칱��J
5��ǆ�>	�0'�?��>�wh��0<i`��?���,ӐE
��S�Cb�'t�ex� ��|).h�}b@�E�[��)p�S�2v:��s�4 �%8�\�'b�*(nLh��� ���1�Jȕy .���F��S��?	3`�#TZ9$ߊo�0��U
�L�<����|�,=C�(^�Q���{�C�u}r��
G�^��Ol��w�ҳ���u׭�@ӥは�0��E��y�0��yJV�A�/�.���o\�~��S3P�l!d�|���ߚclu#�푼9����'��Q�!�dJ�D(H���κa]j�J�e\����tƶ��刋;)��x���88	y�R�H7����#T��0?�Q�����#K�q�n]�T�У3��|pt��Y5�B�+?���r`
�kŰ��FZ���hOX�-��,ȲK�qܧn����s����� *.�Ht��J H����'��dw�x!�	�<���%��L3'�8}���S�R|�x�D�K�ZH4�!�A`ӜYRDmT�C�K�(m�2��OBaĊV�W��q
�(�4��kE3-����2kר|��	�iR�ia)�M
a��o̓^�L���d�x���
O�a�A(����9��Ϟ:|K�i3��I9m4�	�O?F�q�� �K,S�4�yD+M(7�<�:�"O�m{��.A���6�_������Or�E��S���O�>)��W�>���OV!#�`3�9!�I� T8N-f���m����^�8k��Ƕxa�yR��	�<4�f�3���:7���O$LҀ��S �b>9�S��{L�3F��H���Ǥ D�\b��یG���{�2
V8@�%��>�E,^�C��I��!*}��i�s�N�q�I�B�`�`\�!�D� ]�����)'��@Ip/�^�@�'L*A�2��+����'����V�7��C�Lw�:����U����������$����l���[�2Q��(�O�8J����Y�D��-_��Ј*��ɚO�蕰g۟l��Ow�T(�k��M���Ӛ\tP���'��CeM� e�Ru���W�9Nvtc�O <�5*R����aJ�"}���9<�M�s�6+Z�Q��[n�<�T�T�T��bV+�{�������ɞ	���ib!C��g�caڨ�@�}��y�&�R5�� G|bl�TU�'��&쌚V���3AD��|Y�;�i�ά�F��9E���I�0|p�P�F�0$t�ƙ�?�W�gm� K
ߓ0�z ����1(��a2��L,��i��� D�*��Cft���Of%�`0Y�"���5bx� ;1�|�D5cz�$�O����T�@ڲ���+�1|��eX��ӠG#Oq��d�8��\Y"�=I�:�#�c�?=$���N�.vxi`���?[$v!��o[�7Ǒ���Z=� ,{���X�p��hF����ƹZe��0�!�d_?K�A9 �	kl<A�H�.1�F	 ->��R�M��s�)2���>F	��Q��Ax�|��"O��ATN�����@ENT��h(5V���7�).~����'2�x�qA
�:��K���-�Ba�	�^ ��"Gl;J��O�=C<8��+\,R��$4�P�`��4p�ΰun�N(����"'�;"y7���eZ�?�T$I2 B�D����B�fda�3�C�blq��'#������$���IP%�����i�h�caȒ*��S�O�B��w��
h�|	������u�m�Q�漐�O�ԙ����z��'�Ǫ�P0������ԏT�<xȣ��X?Q>�Ӻ�&��H'"a⑦B.����j]|�<�g�	�� �4I&�N� E&Y~}"ဥM0$�(�h��7jǞQ�شl���Ė8;�C�I�(��e]�U��$��"�#Êm�O6�q �DL�'>c�h��-�T�`D
�uXl �b�3�O�a�vI��x�x����Z�&3\�Pcb�0msf��Giǻ��?Q���-_鞅xb���"�1�fm}�lD4|ؤO��5N؋ f�I~����7x-�0���H~NU��p8��)�\ĺ!o���A$8v���Y.�UPr�\��cv�O�u������>E�@af�ZR�T�a��A��Ŭ�O������L���j��n"@�)�_�0 ���ǀ,0x�'�0up �\d��O����1<*��s
�:3��MQLX�5�#�ڑ��)�'�uWC�t;J���D��
k��0��uh��$��2"�& �(Go�:n����
y�h�AA��t���v�>ٴ�"����0G��M�\��t�:W^ؚ�G6�Oԭ"PB8�|��r"ӱX[l�&�ZH����fL�!�ą�x��	�`a�*y(4x���
�s��T)N�!��;���IS^�!�jJ�biP�A�T�X�B�	�-����Viɉ3T(䉒��]`����ϝh���c�>E��'��|9�%�L����z.P�q�'�p�JUI04��I��;h��-Z�'�0s)\�w�����ɏKU��Af�$i��*"�Z,0����� h��x���r���r"�ؖ&9��rG�ݻO��@I�"O�h׮<m
D�טI�Ԁk&�im�!��k�O�\X�[p"dT���6})�I��'G�X�Tǒ����c˳ܒXI�'0�Cg���(M�]�Ǩܿ`n*��'�(��uHJ1pd�� d�(%s�'����@�:���V
�b��<H�'���a�5M��)�F�J*Zs����'$LY���@�I�&�Rv��K���'���؝\�1!�o�U�t=��'��%xFeS� �m+�C]*~�.DJ�'a��Q�*�qs%�Ӿi-l��
�'�ֈ�`/ٻm�(C�aG�SY�	��'��$����Jj�(�`"_�ߨu�'R��%��T����K��d+�R�'�R=#�K	�u��A��Ƌ�,徜��'�F��#��dO���nH�tP�r�'-��2��A=���jw�4w:E!�'�L]��� �5�8PĐ\^n�;
�'��)��LD68�ur)߀Zr�z	�'�
��R�M(}��9p箛^�����'ĬdQ*=o���j5�S�U�6��'#�)���"l(���FI2���'�p�q�)j��AB4l4B钵#�'�:�����SZ��ad'��a �	�'��\31���$�_���	�'O����h�I�L�E�ߥG������ ���a��S��]�rh�Dz���&"ON��3GɆ?9��Y��4j�U��"O�Y�$� `W��Ef��:rf�2�"ON`�т��;��2�I�+m��b��ɕ"FE�#���`���"&��ACP�ą��0Tz&bF�+M�t�p�m:!���~�
�Y��C>|�X� 0%W4!�!�ح @�i�Ь rݮi{�ÃV�!��߲(�0LC�d��2lp䪊�(�!�Dׂ`����@��@�霗��x"K��-M�OⰓ1�	r�D�`'��Uc��cN����$��s�O�fh����8Fdi)�(�1z��M&�ʍ1x��\w�D=D��ϓ�W�r���CZ��<A�2�2n���4Z8z}� E��dݑ?�q5HГ#3�]�t�©��	�O+Le�&h�#2�Y��4SH��K�I�)Lщ�yJ|
��S'����%ݑ�~尅jG-@)>q�'���ǭT:h��iԪ=L�p�)9<�GeW��D����g1򘺁ぃ~Ut����O�|���鋠g�,x� N�� =(e�����r�� £��0|���:9 �f�
9������"+�P �Ӄbjԩȁ�]���)F�Tޟ��цޟɆ���'�'o��1�l����L�:|}���b����O����� 0(��8�C�դ
�R1�Q蘺y���h�3:EXI��U���?��6 �B�:�����A� �5asCC N 6���ɏ��1�� &ml�0E�S��-��$ ������B:�!(	�eܰLC�
�m^�l9�!馜�dbh��'a�	��KH�!�e��Ƣ���۠�bM��'j�8�6���`#M��>[��a$	=w8a�w �6�F�I�#Hꝰ�)S>�0|� FQ#,��{�΅z\�A�蕦�~b��(v,���
M�F�6���4�P��-Bv.��Fמj�v��
��A Ӟ|��iF�eZjI���U7JƦ� CJX�՛�l�)P�b�"�7�UV	��ᤏ��*�H!�t���x�Z�P��~��\I�p�� ӧ/a�qbDKQ�<I��5Z��D)3��9;0�`�Vh�<ـ�،~7&����`0*�K,D�@S5��5>Ɫ7̚ZQ6`�7,8D�qf�,S�q����>z\h�r�6D���sj.S�豈!��;[IX���5D���F�:��覩ؾM΂$h�&7D� (f�ǅ5�
Qa��J~xh:2�6D�T���@ZqS�G�
u��;`$'D��:�0vZp�a��7I��-�M)D�<Pԡ�n���:�:���z�!D��
����mL����uz�����>D�Xpsg�4p��肌6�Q��:D���i�L�n���%I���Aw�"D�|�t��;"c�Q��:�n�J�!D�����>9s&��`�9}�r>D�lB���V<@g�9)��yb�:D��c4�Ge_f=ar��mKҕц)8D�P����JKܥJ�`\h��z�C5D�,�T析nh$���ŗ>���s�>D���sI^�I��ZtbB�ux�+tg;D�p�b�!E*�$@�A>=Т�:D���e��L�%��
�N|:�E9D�$ٶ�<&����	��Ng|<ѲC9D��B�%F�`�fe] y0=R�h!D��*󌂍��׆z�h�"w	-D�YF�3}\�ۆ+{^Ti�Q�&D��H�*Y׀+!�3Q<��#D�|q��¥Dն�z/��:��hU)#D��a� ��B�B��dNԣ�|��#D���/�o7Qb�F���a�� D�$�7O��D������M��Bf!D�Бg�Z[�x��Ɂdʹ�ң=D�xR�HƧC�J��K�C�>�J�.=D�$kK��ୈg� 4>^ �1Q�&D�� � ۺk��Z���m%���QJ%D�(�f/2*��m3'Kh�fI�"�!D�� b�k�Ú3\��"g�G���j�"O� e��[횐
#�K<8���"OIY!⛚[K.1#'��)1�ԣC"O~p��B8Q�R���Ǟ��]�""O�0�5�)P p�;Vf�0��)�"O��iQ�:� ��$%��P4
Hi&"O��ڥ�-Kʙ�b��y�9�"O���J���	1���!E"Oy��mӊ6aTY`� �,� Tk�"O���H��CĈ0"C��,��q��"O��B�M�C%f�qb�ʜ]��u�"O�]j�gU�$��(�|W�h�<IF,R/&��%+ַ��u�p��O�<a� U��A+�|������W�<S�@KF%����%[�(f*�O�<�i�
0`�ϑ(~�!���q�<�P�4����׈ClL���CY�<1!�H>Kt>Ei���s�2q��DS�<a� C
W:^�s��х_���g,H�<y��D�.�()Q���p;HS�H�O�<�`�F�Xވ��g�;2�<��E��H�<р�ۑQ�U8���@�qzsPK�<Ih�N�`��Q,^
��#�$�o�<a��2�|h*E�S�{Z0R��F�<I�����d` �"R�ƹ�Yb�C�I�Z�
�B�f�=^��6S7�C�Y�6��@�^M!a'LLV�C�	
�e�sK�?U�J�F��B�I��D<���U���0!�@� ��C�X�l	H��Ґmf=;��͇d!�䕒5Y�p$`΍ W��+���i^!�J�)~��'b��A���@pS#$R!��
�>�rumN�y�����uR!�$W�7-�p�O�1_�`�4,��83!�d�#S�mj��\��0�'L�r!���"(!�(�"h�[�B`!�ğ�c�bE{bJM`����r��1�!�䑹\�\�Y�N�c���8����!�$
�A��"!ls���b\�!�d�h�F��t�͡�T�CSo0p�!�$�J�r��Kذ\��͕��!��]�H4���$�U68�B���ٓ4�!��N�j��RV�8%
�+p�*E�!��4F{��a�iE�Iڔt�).�!�Z?y�Z��r�D�P#&�[�!�I4].!rP�F2��BԤ��O*!�$ a
��q`lL�z1䌂���*E�!�$�m�����ȺOXU�/5 �!򤊰u�P�iu��[������L&=!��}P���Mƃ!��l���s�!��^9F��V�\'�B+Lvc!��&+���*U5� �z�i�@�!�_�7&e�6%�Z���*Q��p�!�f)�K�s'X��w�D�LX�a�'��	�c��U�]�uW�05~!8�'.j2�ܽ���%��'Y��
�'*��3AJҏ�r��Q���ڔb�'a>�j� :�,T��M�8%
�'k�xk�N}0�׳&�d�' t��7��C9�A��(V�1��'�(�fX����O�Xv*��'zE����,LS����ЖJ0b���'�p�����hL���h	C���p�'��-zg��bEqA�E-Q��<��� �p��	X�HЪ��>V�4QP"Ole D�#6�N�
�"�!Cx����"O
� b
͒t�<�&��g���"OX����x�.L��&X'A�	��"ODd�S�&K86�١78�p���"O������-_��#�l��=İ��"Oʬán�St;��*�B-�"O-�j�!�d$"�E�'�`*@"O� ؅恫S�~8��FU'"�Ac"O��2�����S�:[%z�"O�(��m�-  �vM�z��m��"O��SN� *7Bj�ʍ}q8e��"Oµ8BjG!d��|�G癲&_���"O��릡��� ���L.rx�0�	!D��à62T,���s�<��U�*D���*��t�4$[2�˥.{x0��>D��*#���k(,�T���Bi\,��*O����9i~�ѣI�
n$�=�'"O�Y�`:J���Y��/���;�"ObP���ҿu�*�1�L�d�5��"OT��L*L�saG��C��91�'�����ze:�J�jR�T� �
�'�ѩ���yo~E9��DQ��r
�'!���癸U���+��N�(
�'�����aL��r�+P@ǁL0Jp��'g.�x�闌H��-��%�F����'���p�(V<>�(���3E;�\��'-���UG 2+C��&��(4D�̱1o�q̈�����2�y�7D�ܰ���c�A��#lt�4�:D� 8P�]j�uA�֏W^�;��8D��1�@	3S��a���CψQ��9D����'�G�az�W�MѪPAr�*D�4�@O��<T�$B� > D�#2j*D���c*�5{:>�����|�^�q�o=D�丠a?� �&X
���P�y��6T�")R�`��L'�Q���P��y��8w��"peB��]vm+�yr!#�4�A�Ƀ�����y�N<����$����):��L-�yb!ɊX�����l��R���y2B� A�AZBBN�u@��i�ܯ�y��~Q����ť#��v	$�yRG�%3N�i���0׈tѕ��y"$.5W��3JL�T3�L;U�ف�y�EK�ֵ��-ʎw H�tM� �y��Έn|����J�Ld� d�^��y�a�Q�X�*�A�4h���&�1�y�ީ$\f��V�D��F-��
��y".P<XR�偷K�0H�{�k��y.˪�b9B���~j �ih���yH$uJ�ٔ	�l�XH��T��y��΢D�d�9V�@�2fpK���y�dǽ�����˛.��9��"�yb�V5iXP.��(Q�������ya��[S�A�4�O��E�S�S��y�l�U�f����Z%.]x�HH��y���!��88R/��"�8@�ϙ�yB@ƈ �Ph����%��x��E���y�`�&��,���1R ��@A�y�ʘ;vP�u�W�E�D颖�$�y�E�u�8��"�;�v1K���y"�H�#抌���B_x�\���>�y"M�]��d�����P��؀�΅�y
� � ��I��G�4�+3��?��4"O�LZ�(6-c:ИÏK�1�D�P"Od1���&�ꙁf�[�`���+D"O��l�0��
��(]4aqp"OD�0��<i���a� �p��DB"Ov  ����kۖ4B��ڨy�]�f"OjM:������"@�g9��ks"O<���� o���ɰ䇕 
.�C�"O��R,�=}�b4��c�� Պ�S"O����$c�}����8y�L���"O^���D�3e��pb Cؒ��d�V"O~!I��L**L!��B�
��*�"O�Q��o �v�ms�� �{Q"O.�F�D:�"��ɜZ����"O��+H�\�Bl�#��&t��"OBJ�	�0b��JGӗS?DȖ"O�����O�e�΅�$&R�DΒ̘�"O�`��F�:8LVY����S��J�"Ol�࢜n-���4�ɐ���q�"O��y��	]ʤ�"�M�Lu��"OΤ�0���Q�  q��s�"O �h H�HV�@�W*M2�l���"O���vB	5m҈����A<AOp1 �"O����.K�_v���Я �K=$I�V"O�tc��AtS��j�$�&*���"O���wn�& �(�uAB�Kf��"OJ���5~��D�$�t1�"O��uMüB���؂'�7p��"Ox�#N��#��Qs�˙#��T "Od����8#���D	ON5E"O<���
-��j���5==t�"O�d�s˓Wi;�b�0wR���"OX�P���0g���gÁ�`	c��'@b���8>�l���m�=[�$�EHQ�f(�����>���(���?�QC���?i��?�l�//P��[�Ν�$5Q�[�Hp���-��)����΁�C#�fx���'�"?�����-yb4RN�*t��e�V�Y�,B!���B��ָi5P�0����OJ��٦�oڂq	��#�hΘn[�dZv���;#�-8/O��d;�	u�'x�x#�ɗ�UW�#�2
O`�&���x1�D�*MQL�Z3"����m�sy2�ך$��6-�O����|j�[$�M���,x�Թ�D`ޟ:]Q��A.Y���'b)��g�\��dҧ��L��KׇSDJ��,�ɅBU!��u	WdR6�3יx"��>0 ��[���
�ds׵i4��G��^���	5�x�U�Ǻ05��`��\� >�OhLC��'��;��5���=��4�e��|�����2+BqOL�D�O����<9�����@-DG8 �e��^�"�ݍD.�xr�tӔ�l`≖]�����h��(Ѐ����
��,G�^����'Jr�'H��D�4�b�'����C�/�8İ�(�!pM�uH�e
OT�}�O�?�,�T"�5>�P�S>)�Kr�I$/�L�8�Z+Y��'����iX4�������~,��lĿ��Ol�, Ji�MD.�=���
�,�����Ӥ�?X��X�&�Oq���'��F�}����27��8bl]�N�ΓO���=,O��`��|$B�F��9eȡJ�>y��iW�6��O�Ho�B���O���r�6��e�M�p��x`��ݱ<���ġ&&i���?���?������O��$��/M�����Q����q͒+qȒ�ӂb��3��y8�C�+��%�'��ON}0���lx��� ���V�VA�V�A�i�w��x 񈑸Z����� 領0�(!�D�����D��A҄�wl�J�S��'��6�JҦ�	vy��'t�Oz�"WlI��J		��2j
���(lO>$����� (�C�擽~MtL�c�b���M���i�剅cC$9`�4�?��4AN)t/Ɗe6&J��'�n�0�'�"̑E���'bb��R�\�(���/5����� �%x���mY4l�����_"u"����V�'�|�2'	�7Z��Zbɒ>�h��T
^7mb�KۍRL�!+u�\2O�ܡ@�E]��O�����'_r�g�>7-_#�X�hd�G�0�˅g����o�<q������O�����-M�X-�Gt-��E� �S�O�,��/	�z�bP���"\��0ƅ�-i�6��<1�.	�&LPIs��?�+�be��� hp胑 fxbVI��;�R�3����ɣG�F�0h�!CJ ���3f���ߟ��'{Q2t���@���7c��)'r@$��R�(�a<�d �F�q�蓣>��`Q��J�1�p��
� ���NO���\���S�f�t��#�x"+�'�?ic�io�7�O�����d��U��M�e��-BF����.�'��'�6�rӪ[ l�
�g �Q��Pk�h���u� O�����?5��0�#gg��q�o\Ey2�|r��� ��   �   c   Ĵ���	��ZpG	 �)G��(3��H��R�
O�ظ2a$?�K&����4,a�6�˝.�*�"��ݏ!d!�e(�?����*s�T�oک�?A�']�ʤ��o�y~�۬HUD��Fo�U�~�(S@K�N�rK<���
faKJ>��{G�1qs��/}�p�r��L"g�\�cɁ�@w�	<]�4-�bL%c.�1Hu��i�+=g�5��M��cȻN���9�+�<#�4@���7q?��!�"c߰
��1ҮRb~���Z�h�#/,	����$�ʰ� ��K�@Ԯ`��"����(�dP�O�4��.ҫ|��+��M/s*�1S�^�̓"$Ѱ"�Q��("�|"k�=�t��R�˦]'R��*D5�yBGU�'��Gx��"�� �v&�M(x���&Z/��"<B#'�B��vۢ��V��T��2�Ď�@�h��O�-{���J<��'��hڧ�B�'\D���g �����M+��,Oe"<��I�=|��)�n�E����QJ�Q�\��>iÅ+�-mF�@ (8���<Ŝ$�&�M*"^�4�'���Dx��a��^9,5Ip�B.T8����X܂��#-�nB�#<����O�Ra�"e��P6�G%'+ �V�X��Ox SK<�$�M���X��& �eX�/�H?A�G;�x� O�Yt�ZF��gГ�׈I$ ��	Ӧub�'&h�qq�R�MkJ?u[�H=�Ԥ�9R�Xs�С$D�I�����H9�I�4�B1� D�I�d�=!�O"�$�pj&�p�fĉw'���OV�N4�ɷ�ϋ{s1OR|�����(O�cd٧F �kL�^�0ȵ"O�TcF	�  �*�!򄄁Yb�Ŋt�׺~����&`���!�dW v�p�(��d�ݟ&"!�Ě�l��W�K�bĀ�����-!��\r��ɷxb����Z�O+t"���dOw��4h "O>�CD��JR�I`����Z�s�"O,0XVj�54�����V!�|���"O�h��O�.��с����� �"OP�!dB���iGb�6 ��!�"OL�ajU<���k	x�JI�"O�����X1^�(R�\�W���Q�In�O'����@d2�8����j�����'&,�Ph�z��3���5�ڴ�J>1�|�����)-n	���G�$�P ��4�R����1cg�,��*�a��kCp�7���V�DA`��7����#"x,�G	�6ɸyd�7q��d�ȓEoPD5�]'B��mY���L�&�܄��<4�V��2,��(��H:#Ȅ�`QP���$�	�l'���[:TJȠ�Ԉ@P�C䉷�~�����=fёB���8�2C�ɸ �����#n���G��P<C��9O��恌m�� �T�_<�,C䉏�.�(% [>Դ�st��1z�@C�ɓ[�Z5�+E��xa�0Z}&�lD{���
BoX�$���6��+.�y�Dt	�C��Eh��A���Py��*z��y��ɋu�Ԍp��F�<u�ݷw�����JD�D��$jB�<�팮q���x��u4�`���F�<��D�6K���d�3\����N�g�<A�ܨ
 ���G05oJ92�A{�Ii���O
h�AP��iX0�!5�L7)�N)
�'V`�aJI;@A�q"ďk����'w�p���>*�H��J���hY�''���E̶	�����)�7|�x��' dz���g<�E��{�8L{
�'0��&ղ��%�눦v�ni2
�'��+bD�
e��b/�$|{X�B	�'����肺+��JЩF��TP8�"O���i�+_z�=��+f�:ahp"O�D"W�ɸe՘���l���1"O]��Ȟ�F�jL�R��7⚰R�"O����d�D������v͠4�4"O��az�"p���� �uQ�"O
�xR�9p������$!?�IP Q��G{��i��<4G�r�0�u��r)��V���RgM�>Cx�Y3 U��M)f�6D�� < `iƵg� �J�f�(�0�"OR��F$կC :TK����	��"O�гc�JE�}�M@�]3���"O:�K��B���I��K
p��Y�"Ox�Yq끽[4��J�iہ%b.��c�$#<O0YRӪM+~!���R,h���X0�=D��q $A4kwl��1U��}c`B�O���hOq�d1��A���4��9 ��u��"O�]�"-ڨ��ir$œO�2i�2"O�r�ślh��Q�A(��`A�"O`�r�JͰ-���rw��$�ܠ"�"Of=x�@�2tW�p3B%W�����/LO\D��D%/w����v�A"O���f�����@�
jvA"O������ߤ��ՍD[�а�"O�h�QC� �Ȩ�B\NQ�x��"O�@�oL����T�X�/N��(q"OL���"ޤݢ��@�3&t�:�"O"PRVD`����/��
�T8U"O�h�&��Xk@��%n֝V�:)jf"O,5��Jʥ#�
NA�IЖ4��"O�m�7BM�>�r+�S���p�"O��PW!9��y۷��l�Й��"O �k�
�d �q�߬2�!"O�E�"��OE�!21�d�$�"O����)=(�fpI6*��^��`ٶ"OR*1�Jv�t²��=Yp�q3�"O�

 �-є=S��A���4��"O0��b��%D��S�R����"O\�xGEN7i
�3����*X�e;T"O>H�'@����*:U~�R�"O���p�C����K�˕L�k�"O�ˣ�Q�f:��@�mL6u�b���"O�Pxt�L"=`�8�K��
2б�d"O`����+�@��jJ��a�"OT��a�7c����cS�o��Pd"O��q�
S��0 �ْ4��+�"Oܙc7 �2P�Q�w�5�2"O(,�'�`��)�c�I r'N�RD"O�`{�D�K� y�5ϓ�v��p""O�5�@<B Ȱ�4�U�N��Hw"Of��"�
 o����l�7�v�7"ON�c��(�ڸ�DE����w"O��� "	�:@ZI �E�(�� ��"O�Xd� dL[V`�,i���"OL����9 �r�B����mF�p�"O�ȳ�KD& �(X����Z�4��C"O�9 l@=a��B�FޘFf����"O<��4n�	a,D+D�G`���"O������-WPY�ޣW���g"Ox �O�"
U�&�D����"O<U�QM�Fa���/��æ"O�Г&눃S.(���o��7�TU�e"OF�q�EC�7��p0�ˏB��@�"O��K�D���������k~�Y��"O��H2M���Q�)�����"O����D�����b�I-h]J��"O��ò��3B�x�ʁ�*�\��r"O4L�4i�(��x�UG�m��5�"OT,j��N�HYthI!�A�Ux\��"O�IxU�B�b���&��a���"O^�k�i��g�\!�!��R����"O�EJT��\쩓�N�E56tj�"O� 6̌�7�6i�qm�!-`tق"O� <�9@"C�G�����]9��"O��d��"�̹��ް"uBu0Q"O�tyS��]?fx�#�3L�"O�E���_tDrX"�6f��!��"O� SB��$���;B o��Ż�"O�kO�pt��.J/�m���"O�)�"�Ma���cn@�eb��q"O�iQg������%(_w��`"OI`���$-�68���Fr��"OH9胋�:;��+�]<Sp�e2`"O�Á��Y�Z̑�©e�T�"O�ɘ��haU��-_(�i��*_\!�d��4,���de�{E`%���F�C]!�d�CQ��ke���G��q!S-ǠNY!�dD!=NJ�Q�$_Ӟ� .���Py�(��s�db%��	w����֫f�<a6e�f��ث��9D&�ġ�χh�<a�̜$S�p0�޷C�|8c1�J�<6Qe ���*ʋ !��
s�ZO�<1��V :��x�,�
Q�^ ���r�<QSjI{)�u�6���q���@cf�j�<�Cxή��)�H���[CM�i�<ёG���Lم��$�T��d�c�<�[���8#�
�l�LxP`�<	�Ӂ5��b����>Ԋ��!�^�<1R�F�Z�A�b�ʏd�0��rj�E�<a���\����EZ��L�Z�nRH�<��4Z�~5J��ߚ+����GA�<ɔ ��^U�<C���m��C���~�<�2B*��d���D:{HDm��J�e�<�����~9�u*�V�]!���c�<�Q혘Lq�=���+{�����c�_�<�aH8��Mq�)S%}\��`���[�<	W�J�b6�ct�ˠ!㈍�lM�<��eW?0��<�tL%%��H���`�<	��x�4L@��"?(�uD�_�<ѷ�Ϭ����JXF��Xcr�U�<�S!A)1*"�a���*-�4�ȓ+A��h@m�pS�4���/�f\��_<��볤��z��ĻF�үz�=�ȓirD���R� �1�M�&��̇�d��iխ�/'�pٱ6C��\V�e�ȓJ\ hj��cB�]A&bP�\�ȓ�����3X���@�j���ȓ����$'�4M@�Dh�kM�fJ5��w�R � �V�K��W%J��|�ȓ5BH!�e�&����[褆�DR� �&M�Rޭؔ�E�j<��n���Q�պ((勔M�6,��m�ȓc�k� �%����9.�F��ȓ>��X��%YiD��EQ�'���ȓ�4�)��Q����W��[�z��ȓbt�t �_|�H9�n]S`jX��*4��&�4*�MX�Ȅ8E�ŅƓ]�
�+���f����S �,�"O��آ�N�,�`��@T�gl��c"OL��O��D��dJÎ��%�	q"O,yp׏�XQ� BR�"7�����"O�|�HF�)v>- �J�=�� "O��w��%c<��uԴE�X=)"O|�*�����
(v*Hy����"O�!R�W�ƥ��o�,0}Ή�%"O8�bVdFe�u���5z4X��"O�U� ��-��H��V$=�2h�$"O� \!�OF4��}	 �d4�s"O$�dStZm��*�j *�t"O�z�e�nR�*&,����"Oj<�&�S�T.ZH���µP�&�)�"O�n�dy�╃h�2�h��P&F!�$�`H�Y1RnO1�d��"
O!򤐤2��y�%.��]RrBI��!��Vusѫ'E�1i|�h�A�|!�@:8Ԁ��
�?13�pٷ� 0\�!�d�T=��ّ��#A�RA�OU!��]�6a���aq�A�%ݰR�!��ǣ]`�Ag�oD�"�@��!��N�T�8�B��KZ|@�EN�.�!�Dڅ+��@���f>�����!�D�	S�(��Y�B��0M�N�!�D�!t�Z\�N��܌�1a�ͬ.z!�D �w.j��nȈQ�d�1}�!�dM�	����¡�,���!�L�n�!�$_$P~�$�fJT�� �'ҹe,!�Ɲ�p  �Pe�����3jm!�O�)B^�R�eԯG���f�I=N�!�$�
[/�)��H 7D ����I�!��d�v�1��83�G$�\�!�d�&�p1k0!_)}Tl�<G!�/\.� S6#�a�t�lT�,=!�N�<����GG�s�ꕴt)!�$�+b��h@�-C8�D�fHV7c2!�d˂Rxu�1�S.q�Nx"�LҽW(!���.�!x�	/#�)�%�ǀ#!���S%��"t͏/$h�g��e%!�I1}�<ܘ�G�f�i)���+(!�B�g*�Z/G�
��M��%�w!�άZ4��jW�o㎴���ߢ!�� �,C��2��Gָd˵��1.�!�D��o�&e����"d���	��T�!�����u��� Ri�l�!�dǦ&q8X86�|u�S鋉hZ!��+M�R]�&���a^���,mF!�d��
�X�ã[�{2��Q ߿5'!�ă�H�H]IT�P8?y�騱H��!�D�:wߔAf�B&4m$LsԦ�L�!�Q��ⱂ�OX�$0`�N�!��*B��:�aƎ[���Q�V?�!�dH%G����6��q޴��`���r�!�� 3q��$��>)�*��21T�!�D�QP^�4&�&&���t@�!��+' P���ܒ5��q�GJ5�!�D�:Y�2�,\��Jl0�i]1#�!�$_�� �#&�s6"ȑ�]�!�Z8eb�X��S?S#���F�N!�DR�)M�y2�IƝl>�9�t�Q>=!��,�M�#��@BL�)�tk�'����Y�dhB�ѫ��ɒ�'I6�����0�mE��*d��'M���LA��aAﲍ9�' `���`*�8���V�?�`q�
�'C@����n�K���2��p
�',lu�ݠ%u@�9`�&��+
�'k $Z�C� "�= G�@���8�	�'�@E
6Fi���3�i���
|B�'*��-	/Ql�0:�뛦B�H�'�|��"�vt��CJ}�h!
�'�DMY�CW�
D�1��qp0�	�'(F�k�o\|yҀ��e�Z���S�? ��BTI�4SNf);���s> �q"O��饴�6���y�@���ʽC�"O�����\?�J��GF
�l6�!F"O6�Qv�Z�`���XteŇ!jőG"ODh���/�m��]�]p��2"O��� ą	Q=}#蒋� 8�"O&<�Ș<*h-�%�
�}�
�9�"OZ+��\�0��MS`�׌%��Y�#"O�D����F
�8ƫ�B&���"O|"��O�w�9p��y�NA#�"OD�
0O�9m�̳gD��Fd.`�"O��@��-���r��xaJ��"Od%���9�R"ӂZ_<��R"Ot��uB�.�I�C/~�᳅"O4u��`E'����a�ij�Q "O�X�-X����3�%]���t"O�s@!�' ;��9f�ފZ|���"O�U�6k+c�rM�R��s=���"O��(p'T�`���Zf�k�d"O�*���d�����k��^%ΩQ"O4��V鐹X�(��F�'~����d"O֘"�H¤4m�"+MA���&"O�l���E� AB�&�V� A�"O�D'�I/���RG�]1���e"O��JF &2d`�炏ӊ���q�<�i��@��U���<�4ĂAL�Q�<yq�\%L���ض�*X��x7��J�<ARI�*��D����$��@���C�<	��Άu ��ۄ-W�$#b����	@�<q[�U�G�d�k��%�4��9���R���V��`���.�ȓ-+V@R!"�6*��8Qs!YW�rM��`r��q$5������6 ���۪5r��v�ӗ�"z}��L#��
F��F�� NW
yv��ȓ`"�9�N�_Z�`�P%>s4 ��u�|WbF 	+���� ۤ��ȓ��X��nS?̔ ��Ir]Ȥ��x���ǎ$���Y䯅km�ȓ0� �Á
�i��Ap���Y)�ȓxP:��ܸ0�bH�u�4I�ԇ�9Ly��@B<�S""�Tb�$��*���F�_�Dذ�c�K4�6��@y�
$�ҳt>�#E�3�4�ȓq�$h &D�m�䌩���~X��ȓ2*0���)�%3��K$��tO�̈́�\�<�"]�x�"Gڐ����N@H�<A�ZR�������U�h�p��@�<! �5N$4�&��6����GL�<A'��1B����AN�GƼm��f�<�`-��򁱗��4��A�o�a�<�d�	-N�yR��>V*�ɧZ�<9�Ą
{�X�ᙂ	�vQ!�@q�<9�H��F� U�sC �=`9Ï�T�<�W*\"_����`�C1�daQ�e�<��� Il	�S�5�tIy��a�<If���5�L�5f^LP��fD�<)�Ü���1T)�d��"��V�<Sn�N"�L�u�ӊg�,�ƨ�Z�<� ��J�Y��Ð�(T�<�d�� ~��1�jĈZ!�m�+I�<ٲLځ<Y��D 9nt0;��L�<A�hB�e��@9G�5[iܙz&�	I�<9nB��V�@��W�1��#DC�<� 2�� ܕQ��L��|�T�`t"OR`!'-W>8���r�O�b͓�"O�����>I h,��.,��4B�"O���a��6A�U���լ{t��"O�y�A��`��0UmW+<^ hI"OTe��M��[p��V6n�L�&"O�a�J�=h`�x��A�0]h�"OZ|S�Y�t^����]�2/���"O*�xX)n"�TlܔX�8(���{�<9�p��%��[*��#�^�<��Dݙ����Uf�i`�Tc�.Oq�<����P���W��	H�ꄆ�f�<ٵfK�S�P9ӀhIGr]�w��\�<�"F�~��L;P�XE$ �#�!�L�<9P	@�|������M9HU�Ad�b�<!!�ua�e�k��٩���`�R��S�P7�Jݔ���ĠbItY��\�ⴊ�!U%�Bܨ���b���@ᤤ���3� ,�d��R���ȓ^	V������8D��I\&:���ȓLv <Z��ڮ,���t�"wn������ ��B9~�8�&*lͪńȓ_'�ɓC/!8�Uȱ��=v.0��ȓ�0|��ɼ+M �#�J?-�����}L!q�@�GF̩����8�ި�ȓ8�5s� =~���%F�p�F̆ȓ�N8c�����Pv�Q��-���@�jE�X�krq����$(Ň��n�1�,"�h��fAB�Jt�ȓ)5�T��I
����m�[�bl�ȓ K�iЖ���U2���4�[�&ŅȓZO�4p)�����1���?F]tP�ȓjZ��t�1|��°�e��9��o"���C�v�4 �-`k�ńȓ'}P��aBF'W>��C��n�,�ȓQ�	�ɉ
{�9yB��g�ɇ�)��,K��V;h� P!��"��|��IRJ��ʎ��� 	o6Z����Hq�)²?.0z��1�)��k�ĠG
_C�h1* �؟
���ȓXx|* ��$W�t��!P�-
u�ȓ`�U�t��%�px�&.4���ȓ%
�بJL;0|~h0�e�*2n��]���J��ÿ���O$�|��ȓW�U����N��{�Nثn,����]g�u`�FC�P���{$O�rWvP�ȓaO����.�}H�����*w��y��^�E�tI>L�iu) 'e^ �ȓ��d�B,&�  	�._24h��T��!VDC#.�k$�'.�&q�ȓ:iJ��kKA��a���j!��ȓ,D ]�	��A9[3+�h��T�ȓ�Vx(��N�TS��2 �X�?��݇ȓS@�ZQk=#��P�	Se���ȓ:�~!�`/ǁ_c����4��7,�ݫRk��as�"�n�s6l��q�8�%Ă�:��=�R��Z�9��{wT��'�:3�@B'C���	�ȓzp���bV$=},�"���P
\�ȓ�^\)�
 f�lJ�(��E�����7Hݩ�� ޙRq�U=h FP��*�m��Qy4|R��ZNT�"O"��7 �d1c��+h��br"O6!�Cj�@�e��T����b"O� �]�`ɚ8E�A���\�����"O:�:�
�B&��s#�P��+�"O�t��&��I���:Ζ�q�"O�=aU�K�a�NR�����*�"O���!��`��FKN�\� q�"O�HR'	�Xn���A�	� Zf"O:I����N��M2EH΋K
UR"OڑI����f䉒��	�P ��"O�����;(�І �
&��"U"O�JQH�rڼP'B��1�|4!`"O0��� L8P��
�p�`$�1"O��x׌�U4" �؞r�:�r�"OX���//��08�l�*$���p�"O^��qa�8mÄ�t�V9��x�"O0�q2�/U^�����\(0��iK "O
��M��P���OQ!�}��"O�y�J�?��г�Ƃ��"O�=�v�Z<L�
F��/W 8qy�"O�!�2�ڽ����)�� M�؋�"Ov ��ˆu��qkaIC38VX���"O�T�G��^���ÓHȼK^n�"ONe[���6`�d�VHTfH�l��"OTcF��.WtI���&WH��"Ox1#$�*j�V%�!� �l8��)�"OX0Q$-�6rP�}�����"OV�hW�˃C�h�'b�<�5�d"O~墄2+���t!�5�L�"Oؐj�ɔ<�6ՠ�<	 �e�D"Of�Y�Dޜd�BP�ӢF�\��1"O0���MxV�|�K�y��R�"O�eY�D<?�Z���g��	LT�"O�E�� ޙ 踱�� ~)�Ē"Oe9�֛+���hΨ0�ԑ�"Om�K�?�R�Y���E.N27"O~�+Ac�,6��f�6ʺՂ"O^�	���7 ���6s�%�W"Od@+�]�g��t��*	>!Ȉ�6"O��DES�-'&���*��]��p`�"O0L�Ё�4��A�TCD�F���"O^e�-ʱ^�}�2c�+{�8B"O�prƃ��&M:p�G��oz`�`"O~�[S��
X��RL��P�"O�䑧q�<$���?a���z6"O<�C[�M��䃶���X-�"O��Ȥ,�U0N�s����%'T��'"O��tHڄ����/
7^	�Q��"OD����ņp)X$:��� bZy�7"O9k�U-B�`cF�������"O��	���NjU�&K5�N�C7"O��X�*�>w4x%���-�
�"OI �J�I�x�h�g�(�Խ��"O�1�g�7^��  �B|�l0"O2Ys�čNO
1�g&�U����"O��+фHV3�DkD���Z
�A"O�<�`gՐR���D؉�\H�"O�څ�,7�Q�-��y�RQ�'"Oִk�,W)���!�m�h��+�"On	� �i���X1�B(x���X�"O�Öh��)�&�|��`�"O�M�Ǉ�榙rD�;k�n��"O��0$̧c $q�)� ���r�"O����$V��1��Ċ�^]�S"Oڈ�ul�k�X�B\
I�L[�"O�Q���W�02j�PW�_� �B"O� �Ŏןr�L1�J�7�t��"O>�����Y�ݺD�^l"O~��ۺ���{�M͒y�>���"O\��KK1X"`b ,�<� �"O�8�S��?Df �1�90oN<�!"O2�2a��9�A��1@p �*D"O�p�� @r ���U���!D"O�(��"ѱGXX r)-:	�T�"O��
��RF�LT���j�2ѣ�"O�0sQ�˳Vx��3�LK1W�Ʊ�P"OFB��bS`ٸ#A�L�<!1�"O`	`B��;!�(�� �]T� ��"O��i�Y��bd��1DP0,;�"ODT0�FK8N�L!� Jݥ*��[�"O\d�ʬP��'H2c����"Or����ʛ��݃R�߯X8| j1"O,�;� �}K��p�FQ�~'�H��"O"m���+w��H��2 �jb"OZ=!�j�Tm�f Jh���s"O��Si��=������Nv��F"O��ki��?�QR�*U��E�"O^�rf�C3De0F��
��ٓow!�$"'�l����,b�4h��@I6A�!�]�K�	��g�
 8tE�)Z{!�D=� ���I�-�
��e\�E�!�D��W}����a_6_L�@��D�+!�$�2AF��D>e�U"wB��!�͜@ ��(��.+.�`v@� !򤎖&�xІm	K��Hy�V5f!��Z1S�萃��J��}( -��!�D�	��!��'�,U�����[�!�>]\�;.��Ih�=C�(Y�Nu!�$P�&n6d�G�.MP����(N)of!�dO.q�
;�ߟxFPa�c�3e{!�݁[m�������*�h��T�[r!�D�H����p��e	�0��Nl!�d��B:��z�ϑ�M�$��1c!��O�3w�l�F�M�7l�XKS� �!��](>��Mt���Qj�0B��^)9�!�d\��MQ�)\L(��$�O!��q�@S�K�}7��3�� ]!��T5#�~ ��%ַ[�����_"G!�d��v$E���R��r���W!���"ߴCô����]8vڀ��ȓ.�Q�덉t��Ї��1-b���;&�	�פY)e��pGO��z4����')�0��N�g�����Y+X�u�ȓ#� �[�Ҏ��'��&[�L��(X��y L�A���HGB�f�Ȅȓt&\:E�"$A��@��]�����}R���A��?���e��f�&l�ȓ%u��`@�ʈN��%�vA($#d�ȓo"� �9D�0�G#F�4ر�ȓJ�x�SmO����Kg�A�:���@E���i���F^�4X���q�l���K<��{�m�1J�����r5�Â�'�J���nG������G�C�S�^���i�$8����)E�p{���cd�}Âl��g�ƍ��~��9Bn�)wG�����7Q���h�"��Eߌ�,1a3o^�;<���z�H�P�N��`��D���M��-?�Q��aJ�ȝ�ቍZ���ȓJf�ɸQ�Sǚ�r1}�����S�? �y���՗dN�=;�+��"�!�e"O�����K{~����I�YFTZ�"OJ�
3��!I�8$Y������
�"Oحa�i��<�0�J�S	 ��"O$��B�7�z��c�&L��S�"OV`3L��vaz�0�	-)ʢ@k�"O�<���C=���Zc��!��й"O�xbl*a
��� �>Mh�"O^�S�eZ.p�h��}	��E"O`��� e�݁2�@%%b�Ix"O��`���FOL@�V<Y���"O��
ˆyF��ѷ �)Lפ���"Olh�o45�̑s�JҐs���"OT�j4�P�H�˜4QR�B�"O � ��E6\�@ݺ��-f.�a�e"O�a�J�?Swn-6
S�&)0�"O�Q9�Y9o�#P�ґH ��"Of�a�.ҦxD<��Ԕn��X�"O4`r�$���`	����'V8�]K"Ox9D���32��"q��<{�N��2"O��"�m�X��%�^c`�Ʒ�yR&�'	�l�Xgӏ1L�#�C���y�o�0X��5�&)���%����:�y�mC7'��C��_�����&�y�F��(�RY*��V�P]S��y���B�,8êHp:�(� ȡ�y��	P��t���]1B�n����y��Lz���Rc(��U<�yRf��]Ռ�J�nƴHp�=�����yB��5����.�X�nu8��U��yb�f�X�xV��|L䕹��A �y2�O'�M�ޤr���aꝊ�yb��"P��{tbO�2��XjVB�y�)B�T�c���/E>��ݖ�y�ʖ(wF��h��'�=�!Ǟ�y�`�q�9q���-� 
!H�<�y�lP-F����m��	$�S�g��y�+֘	 �4�GJV�ܱ(��y�Θ�S��Q�.I  /V��y�-��>5���9�����Ƅ��y2��<c�tBV�Ј=��q3E�Ҽ�y�)�z�^}1��G4�N�JT"�.�yaC$
�j��0�33G%S�0�y"�T}d�͋>\\��"֢�yB��5F"ų�`> M~̊�	!�y��V���dTn�8̘��#�y���QP��2BJc��Xdl��y���"S�q��E�C�ʙ�#(X�y"-�_��}b` S{|���X?�y�E5� ��	&N讈�v���y*�M��DX�o�AE�e �/�y�E�J	9��&ݨ�b�(�y�C9V�@m "��	*<\ԁU2�y޼'�qyF��Y<9S�R��yb�ΟlR�]1�Lq��K2���yb�Egm�(���\ VD��1�ٝ�y��6EVfl����&����Y��y��?����$�fn��Qk��y"EP�H`x�:��؀{��<iQCC�yi�+�(�2ĊC�s8ء`�G�4�yRψ�.�(Q���\�g�p�ʕK���yBnU�#.�Q���ūW�*��E��y͞"p�
��i Z�=��(�y��5S��v�̗G���q4b���y
� (d��d�-^x�Ő�j�:G�����"O���`M�b���ʠ� �yuP騴"O����a`�	C�\���"O��a�B1>l<���ܙcv�� �"O�AY�C(����H�|9L�z!"O�̊��9nh��RV>{n�[R"O!:Tc[solx��5�@�X�"Op5y.E�:4��o��R��0ȃ"O��d��9��ǆ�Ev�q�"Ob�8 "Ʋ<t�z�g�c��L��"O   ����I"ڴ�ԦJ�gЙy�"O�U��'�8P�t�aE���l�i'"O��2T!0^�r�q��h���"O,��n@
a n8b�Ɠc򀐐q"O ����R ��G��34�0c�"O�̓�CA8a���ȣ �+���V"OHEj2��
%l�Ȁ�� 8� ���"Oj��Cf�+wĎ�  L3d��@u"OZ�#�d� 	���U8:ap}q�"OZ4�k�0?4)���#N~��q"OB��1M׭s#8�qƠ�Y��A&"O�İAT�D44�Jc�[
�ܨ�0"O�P��mC
\�V��a��u�V��"O�(׌�%��Z`�.I̼�JE"O<�
��~�
As$	
8F����"O�9)a�ƩKID ���پG9�d�!"O���C�H�Q$�@i2�	��"O
Hd.N4[1�8��,��!V@�"O��8���p��s����usz��"O�X���8e�Б�o�	D8F�K$"O��� �W=r6�� a�0=ҽС"O��HF@X8Q���&{-���"O��Xe�ի*�@dSԄ/J�p"O��Ye	�p�B�3uDܓJq����"OPYvH�9c8�ܪ%B3k�L 1"O�H�O�d*�q��D¶n�a"O�H���N��2�dЧ:�d�"�"O�	��$��-�TX��DY�b2��"O���F�y��9��׌o�\�00"O,�����0���B�ۈ0���{U"O�d�����4����N$����"O�R��P��p���]8��7"O�}�$�F�$p~�a��#i�YA7"O�!��j� KPYTJ 4 ���!"OXa�.J8r`P!iّ/C
��V"O�x��
���Ia(ɡL�=x"O4��&4BzGh�RD��6"O�dD�
2Xb(��-�)ta��"O*�a�nx\��Bm23-��"O�Lj���� �	a2暬C�`�"Ob�c��ұP�J��q�ƨV&�Y�D"O�-�o? q��?2H�Z�"O�䋧��6Ʉ�I��@L~��@"O���*DK*�q�`֨^i �W"O��'��o�6��A�<mg2Q
T"OtP�!-[&R�踈��[�C�Ƅ��"O�i��KU�<h��Qp�;,�Rx��"O1cag �z�~�#�,�9x���4"O�� dDV?$��&�]|���"O�D��
�<a�䢠B��6R~|�"O ̫׆F�RP25�ک�F)�G"O@p��2�8��wc	6u䤂c"O,���I�'J��$b��J�mdl�0"O4%��`����k��w�x��"O� @y��Ђ#��X �K�.� ��"O��c�D����!��/��I'"O�%���B�[��8�N�(�E�g"O���r��6e:칃��4>�L*a"O�Q;��	 s�Dx���MM3Jx�%"O<ի3��!f҄xW<=(<�Ҧ"OT��d� &A�Q���X�7Ф"O�HAtNԊ?Q�� %N%Nz Z�"Oޥ8��/:�����ޮ+5�Y�"O�-`֎Q�����F՞(��-�!"O�c�I�$w�`H�#�A�N��hh@"Oz<J��Ճ�m@����e��h�"O���UA�E��G��X�h"�"O�=��@ޗ3�Q�늬	��K�"O�g�Ї*�e��)c}���#"O0��� �o¸	�%ȇ�2E(͠�"OP5
2苊"4�����[�Z%r�"OTM�e�\�u$�1�g`͝��9�"O��x�'&�$#�¯����g"OB�#�-F�J�i�nY�d��ᙅ"O�Y��m�K*�!��0d��P8�"O�p��V/GMP�"�ތZ"O���ծ�<�(G
���`0R"Oި�% J�v�҅b�,�o��u��"O�����ўK�$P��[�C��ݚ�"OP��&�scb� �+q��U"O��� �ƘgD�J��$��b"O����L4@�2����Wuz0�W"O�(�r��>w�V��B���Ao�8��"O�1	�f5�l��ċ&P���"Oz[�!��s�t`c!)[ް)��"O��bsŌ�h���胬��є"O ���q�;���	'�h�&"O`8r�D��G��b%o:!��I!�"O���π.)�0�#�-'9���p�"OL��  �?� !�P�9�9"O�1A���?}���Ѭ˗!�L j�"O�I��-�� ɛ�k/�j2�"O�|��[�G"
��R����"Oy�bF�P՞�U�PUI�V"O�\ ��A(K�2Xpc�f�XK�"Oִbe�>o�4M�$�֐?� �f"ONp3�@1g�~�KE腼���1!�N�	V=�`Ɩ�H� eXc+��Y#!�Ħ�(pG@}Bl �T'[e!���,{��	�a�qs�J���Z!�$۞g��@ۂF�@��I8T&#@!�d�#F:B��a�w��k&P�r[!�$�25"��'F��zi��ER�!��<���	6�
� rt�E+y�!��̥co��A�i+G�k���2�!��ܬX�8
��ɜE<||ꑈ�[U�'�D��I�t�(E �MU.P��cʱ��B��Lp�5+�4Z~�s&��;	��'�ў�?)�2�M�+����,�8nH �R��:D�����I7v� p"K[5c��`fC�>��)ҧ2�h'�(]�@��9^�����m�~��-	� }�Yc�HY����%�h��I�m{���hB0x�.ٙ�ֆ����D#ғ[5~�9�GA3Hw�d�P+?`D�Ɠ�6�#��iB�뇫_�LH��	�'E�q+�1{��
$��K���(�'�P���ɇ`n���"@�6ي�'�pպ�
$P�v�Z�Z�%�f���� >��� Q�$�&Mj��^�O-(�B�"O4��`i�.�V��Jίk�,PE"O�9@� ׏p2����i�{�А�"O�%���Ǡ~�ҩ��G���>��{"�I�4Hdh��>'{؁�Hͯ�*݆�	I�I�jЌ(��7L�m����zF��hO�>�*�mG�1�h�.2�R���b3D�(�f�Z6%���*�9p��q(=D�\ȓ'_X���C"T�M �z�7�O�9��|7�����Ea�AJ�)�ql����ēdF�#>�'�H�jˏ`St�q��U,~v�,Ӊy\����[��<��kH�&�<h���[]}(fę+�0<Y��ʽ�$��'�#@��ҥ��-IvB6�7������X�'���ꇋH4�"`
�lJ�Pl0�'� ��բşoy}��mΟq�n��
�'
v���"S��.Ukb��2pE�	j�{��)�	@��w�˴:�`<(%l�<F��a�:����w��v+��1� �!�'��'C��r���O
ͫ���V:,�����'�jXC���;6��իGC^�cNv�X��$���Й���H���hr����-�Ş_�����<-�])S̬8O.��Y��(�'�]��n�6�\"�>�E~��d.B�o�Pp�n]��P�H$�[�<���C�7��q���;=j�PdFQ�'1� �O�T�rf�fm"�ڻ}�Ѐ��'Y�M���A�L4Cm�|J�)�A�iZ�"~Γ��ɓ���Y`<� �J�d�6Y�?���~R1�\�UD9�ڄUSt9�ÁX}R�'��5S����jp�ȅ$� � 
�'I�����_*�z��>O
�+�'~49�6�ӂ�H�Y�BZ����1�Y��%�2&抺D^M��"O����&�*o7"\�$e֐��p:q�i��)�禵R��:4#2�SR�˅j�~`臃'D��8$�E�@f��V̈�hlBR��>ɳOc��=�}���V�d�`�)؏Q[~�0U'S8��IZ}���"5�\�@�B�����(��yL�R��cU���|�j�OL.�y2����њt��
B�4᷀��p>iN<�2�A;EĪ�:�'� f��+��Y�<a"EX�k"��q���}J�ysV#�j�'@ўʧ���r#λ9J\��?�H���'铮?E��'D���K�T���bmRNdFP
�'I|D�Ũ�,�4ZW��A�f���D&,O�,ӕ�
 {���Mo�!���'��'���M_4n�|r`aD�}Dj��*/$��)�DJ�&�̍�ć���*q�`.*y��<�O�@�
+���bg+�I�X�9�'Z�y��hZ�cj^��ٵ,\����y��)�S0��ɳ��9�p�
᫇� ��"<	�>�S��i�Ǌ��_6k:M�r"�!!��B䉷]<��ԄV�� ���@B�by[������ۈ���Z5K�,�xM��%o��}Q���Jyb���y�6�4	Z1Pu���t�ʰD���y��u��$Ţ-��xp���X�RXꔄ�{������Ex��	�21(�3%��>�:D{���,�1O���,��'�'3B"gCK'��-�4g�q�'Ŗ�We<���!�oվ'�����'����C�����'$*��4�Px���29v-��MY`&���b\�M[���'��|Rc$�7D���G�"��	b�'"���B3(��c'��|}z�'o�S(�%J��u*���t��O��=E�� ���1�]�=~�dۡ|bMpr"On��㎝�l��������R���"O�ERa���Ī��F�5�*t�`�Zj�8�'�إ!��V���x���f*B�J�'!ў�I�@M�"N�r�EI\@���*�d�7��'q�d��N{�	�e��<�4|c%�&�O07��<��Gα��=)E�
�y�p�hIC?)�Ox��N?Ɍ��'�X�P��+��&F�$x��،��|�Ԣ~R�/�`�X�gɚ�g�n����N[�<)�,*J,�jvQpvԸ"�o��P��I�<�.E�6����#��<I�d"P�h�������:'�"ŉ����Y�+
��!�dY5)#jy���)n����D��<Yy�\�W�)
B������� �M���H�O	a�<�%G�n^�jpC�00B�1���s�<y@���}��`aLH�M�T8d��f�<nȘk@m����&'����u��|�<��CO�>������a2B��DǔA�<iP#�)xP�\4��c4�a�V�<��
?/�e��G�9OY�)��HU�<95Nܷ! H��DH��]�A��jR�<���_�xۂ�ƳQ�<����I�<9�-+op!�e�
p�𻐎@�<a�jW�@�j|a�O,	蔘k��x�<�F�E ��Q���#����r�<��B�H��<�A��#$քQ:"�o�<�S��'[P�s��æDq3��(D�\)��$<d� �/��"�%D���M֕8��#=`��AA(D�XQ*C�[�����O%Mh�9�D`$D�|�q�95v�#�B[�k��6D�b�ɓ�A�Jm���2��8�K7D����ʷY&�Y1*	���[&h3D��mM�N���1OF�7�����3D���E����R5�qq8P�F0D�`�L�*Έ�6c@"C�,仃(#D���BG�^�y������{�mn����*N�9��N(�u�T�^���'������n��\�	�����'e�9y�%Ԍ,�(Xl��Q�ݴ��'�l�)�3}���x=���m=f��2W~؟<�����c�Y�i��d)a��q͘�s�OZ�i��;X��@O��C"�x[��'��O�p�ƍ�/s*p ʲ��$6F�;�"O��*��T`h8���!�v��A�"O"�i�mTu�-���T�m�Ι{v"Olm�A�5r��tã�Ŋ5H��"OvY��F'1V��E�T8/���i��'�Ě9�| �ʌb5�}�#'�N!��N�~Ò` 	�% ((�p윴A=!��3=� ( F�N��J��#!��?p.�:V/���Ѡ(O�!!�$(:2`;ӌ���hXrR��T�!��:�,���7k���%�cH!�O?�zM#fM+.���I�k0!�/�,i��Ǻ��d!�C�:)!�P8k�EYT��=��L�$��X!!�E7H��q�G�-%�������'!�D�#9�[��ܠK4X��OE��!�dɣsP��A*Z�oT��aϸr�!�R$6"��cd�]&�=2��C?���_3������ ~5��:p%���y�Ð�k�F��o��s="-y�Nȇ�y"��"ܖ8�aɁ]���ֆE��y
� ��fb�0i|N!�dԮ`�5SE"O*����y�b�r���8��l��"O�LЩ{�ݒ7
@�h�8s"O~`8�h�2F��"%"����E�b"O��H%Dɬ5Y`�Kp�I/a�$�Z�"O���IK�n`�AS4O��~ZE� "O>�3� @�zE�V���G����A"O�hs�o^'�D��Ԭ��B�&!�&"O̼8��
�����d�<��"O�����S�+/�4X�-G3n�U�t"O�Da��2c�"�P78�f��"O<݀�Ҁ(�|-CL�}5(T�%"OdÁ��4��F��<b�d�S0"O*��Ui�*��8c2�1����"OXM�AE�wp
���g8���!�"Odl�t��1"
�ؔL��h��\E"OL��g�E�F�i �ղt�����"O�\ر��7l2�lc��>� �5"O��¶"��c�*���Ź.��)�"OjH
�S�rՔ��5řn-��"O��K����� �3d\�Q*��y�"OX�S�Gׂ����6�Ǆ���!S"O89��,)3N�m�����"O�г�N[/=���R�F��jJ`"O���iM�Q��m�2�Ni�Bm��"O>�Ad#R�V�p�pbWW6D�ٱB�C9<���' �`��b$\�5nc;�z�rT�!D�@夑�G�B,�2%��,�$@��-:D�к`,Ŧ_���'E��0�`5,D�`�._#!Ϯ�w���܋��*D��歛�FW��w��q��Dy%*O&a������k3�ż _f���"O��&�ZX
���Z0�2"O��!`�B�P���F�Q2w�$y#�"O2<�g疢efzx�d4V�Zy��"O҉��ˁ�;r	*$ܝ��"O�S(#-�H��O�6�@4�"OR���@=�.�<x�JX�"O��Rb� Q,�m��#5]F.�4"O6�)$%�q�d ���ߎ/>|�"ON��Tg�L�Zr��RPaȑ"O�3W⊭rfE@F��9�,u�"O��;rNܺI�\L�b^�f��p�"O
�6�ėB� ����s���3�"Ope`��%��H�1)Ҥ� ��D"OH�)��K�P��|�ዕ�v�8H��"O`�X�K N���hP(0Ūp��'� ���$�9.�ɧ��z	v`Q�SP�O�|�T�d�;D���R�2|H��P�є5�J����>�cJ����At"$<O�$�4!QHT��ic����'Q��!�ό�*N(Y���t���+Ұw8T1�P�*!�D�/^��EJ��BP��8�Q�X�3L*J��%ʒR�'}�\��gP9 �t����� K*��ȓS��J�{G4=��I�:�L�:ş�Q4XѷL��)�矜K�nK�iN����،pD�x M3D���s��?i�59?h�ҥB77��	4Y�8����Ǔ+����I%FNH��ែ=^�Q���h������XֺAc�	�\~%ffK�^e��yc
�b*h�B��7$��#KV2��tӂb!%r,�0�h"�"�*�K��0��dÊ�de\y�DD��	������y"LA�H�|j3�	@��dإ�Ֆ ��4&5���(T�<E��8��*�ǒ<'p�|��a�d�0%�ȓ3]� �!f\�J�m�� ��U�\i�'��E���=����!��pGF �$5)Cʆ�KT����JP5 2�*� ���T��(��)5
̟A/&�h��'��bP*�S�a|A� &(�g��[_����T#��=q@k˹=e^�J'�Oy��,#f��I����r"O<8S4jU�,� e\�l�ބj����6FiL���!#S��"}ҐK�:�"�yv)M�m\�P�7i�b��Қ/ټh�O2���հn��e)T@�9���c�"L�H%�f(ٔFL�'�8IG�,O�`Q"n ��e@�G�g|P�6g����Y�2��.�3�� H�z���}`���&b�.\��M��l<2����.�p<�ҵj�� ȸH�|U��	�q�<�Ѧ�)}�������""��z�M�3h�6���x=���)5掑CUΑ>u�џ�hÒ*���{&��y��ۮyR�����ҥcWh��̸'�ح{t�@��b��铧|��|�B선&�J�X�ܘ+��ʓ���J���ui�D�
ç|�p]#��)�l�I���7NV7�p	��Z�`xS�<1��D'cĚP��+G�n?��!�m�&@|�'���p�fI4"?�ϸ'� s��&V�0#C��^�D���n��%��q�E��0h�<C�V_�@�����#�p�sAH()���Â�� `%��*���<�����D�xDց�?�E(�	w�����	��6�t��T��A�]#:AZ&�V�:%�ݺ�f�%]��$�5�?�F͖�=��@�R�0r�F���<���4f�+���m�OX4T 1�ٕ<N�=�'.؁��t(楃���E��Z����O��(��| �'2td��e�$�P��Үj5Jm�'LM�C�4Tɒh �.g��i���%;�e5l�Sdj�Z�Oڗ\H]F}��Ц0T�ҟ%Y�Ȕ&
�O�LP�jS!��Ē&SŨT���V�
e����"�(Ā`��B�EAҎD{�8��"�Oti�t�1���G�[g�������H��� ��O�,sU,�/+�,y��'�ּ�6�/����LL4D��CV_N�<�DG\}Ӵ�k%%Ȳ6��|(��Ox�홗��WV�$c�'�d��qw�U�vNU�����#@6w�4cC�y�t܄�	�dj���	BGTz�jU��YD�Jw�$t�1qeᆨS�.���=lO����νu1��0�*N-��D�b����9���G���yb���;���c�ʬx?���*Ѥ���@إ��.!G�4q�' $i8'_�ItZ=���� �$�v�$|��d�On�����<�����{ޭZ�ؾRT�4���\�,p\#l6D���&W�.^����^�\��� ym|�Ƀ9��u�'���/W�$Ex2�ؘUJ��
�\?\�Z89"��ϰ=�ǋW	"-Td�)�OVu�׌B�� �0D�öU
�)2v"ON5gS�*���C�8

ɢ��@��`����h���2�� 8a�����}����"O8q���$:*&]/)�I	G��=_�}pP�OxAq����yჅ��?:6f�/(��T5��-j�E�Q1.�kd��5aĄx�"O	b���N��Z�%�&���;Ph�!4ˢ�ؔ �O�`
����O��R�O�� �wc��h�#
A����!��p�Ĉh�'�f�CŖ.ij� �����P e�ր8Vf����,�҉A�NE#R!b�3%Vo�'��`���"$����Y,w`��;	�%����3�X.th��k��
}9�ف���x�"���?M|Pу����i2�Olt[�˘�Z�)ӷ�C[T`I��|��WLP�G�#���3�E]3xW"t���V��oԾJ�R2���%��%*�g
��y�oӘG	��Xf��=�jɹQ�ʦ2�.�A4�]�cl��#pL�?�lr�/3�SR"�ͻo�c�H��NWLm��Q�w_���Ɠa��|y��5\Hأe=���tn��x�e�>\<N���,L��T0A)�We�,yE�!��u�Ƭ�ƸЅ�I#��]�f�U̬�15&O�F����C>6�jRDR=6<�I���D�(�C��'\̔���L�F<m�C���}��4�O>�c+~��,�%��Y��l1@dS�:�f���H�~�YYF��2�&����7u�<��ȟ�#y
���ݒ,�@�G�_�K��a��M�-�ͥz�������F�p�X�]_d�r��u��8��L�?R�B��/��5)a��J��xB�ٕh�H�GG`��.Kx8)��ʍ4@ ݳ�M����O�Șg�^0G�5� F̼StL]97�'��v�5�F��'����Gi��`���L���Y���'� ����86�|42C����fΧW.�'9��c�̟J6�T���G�f����[9`9���O9���+ r��i��O5b�
���'餩aA�Px�f��5]Z��2��5�)� Wj��d����>��O������<�B�'=�иB���i`�@��BHM(<�&"�EVb�sХS>$�h�q�#�L�X��嗽X>�k�n�t;��tDCZz#>���0���5����6�A�	S8�ȸ��W&C8f󔇅'PFlP��� ����n�����B ��#~~L��#���BŁ1�'tzVb	/R/Nh��Es�H���F�߹3�� 0��C�F�R�5��
k���+��?E �+W}6	����;�Z�q�M!D����Z� �ȕ��(@?^5�)��o*�E0���Y��PEP� �b?}A�����y"C�8��H��L߁ ��T)�����xGT�j#�y��k×�$�1�O^�L��V�n�"`)A�ff�Hٵ�
h$Q���fb��y�xy�Ҧ 펽��&R,!�򰊇��Q�'��k6���M����c*��W�`������s'�kĚ�Yu�V}{"�<ٗ��
��S/,}�.�)N4�����.j�扊�ۈ��'�N�X3��s&Bm��_�9�rY#%��tbN���0R���4����$�Tfz\xblR%l|���)�'�$U*��.nѸ���'\��*HӤ rɑ��v��X��<I�HO�>]\�£%D� I �lS�`��\�'R��AͰH��ϸ'Tj����<0޽�3���-�F��{����cC]�;�4�A���Z�d���S�Щ��h�R��D��M��fY<;	�a�,�Z~�4
��½�~����e���y��3 �:OL��O����g�X�t���<��.P������\�8s��B �Sg�Z
�|�T�=���P���#l	�L1�Ác��5�'��9��EA��!���O]fH1c흿?��hg��|E+O��փI��=�` ��+�t �/��U!��JP� З',^�x�)D���M3�łS��i  ����|9�`�V�:4&�sqdB�v#b��*�r�br���e�d*���"�R�B5N�%��0sVn�<AUK�d���z�����c?)8W��}5���-^�^� V�7O���*�`�RN�\Z' (\D�3 ���q&,%t���`�>��eP�'�f#}�'N�l��B�1h ��k��a>�d�N��PB-W$*�x%��?����AOA��7D� �2$Bc�<0h������� `#W�& B���Ғ�a�`˃ �`q� �(�z�Ĉ,]�4��) p\e�ˌ7�>L�QGK?��t���۾SE�Ȅ��|F�	��@8�pAhB@Ԩ,h���=1�7���cr�:`Υ��K"�S�El	���5|_NL	R��	p8B�	*
�@m�a�*s:��LD�����P*U�=��GÑm�@��j?�'��V^��!5@[?+ �းO�!�[9V�tS0��+P�`��b�d�1�L�9<�b�oǟ+�]`6�;�����鐏<�@���HO�:B��	X�������ʞ�W���hf��8f5D��!�3K^]#��dr΍����<j�K�f<9>�����o/�c���Agєk%��I1cG>fFݻ���i�ӕ2i�a0geƬ.� ��7�C�l&B�I&L��y�vÒ�|��	���M"Pz�y�4�j96	��\!-��$�'>�'�򄝫aNZ�[��	�j��$�2�!�$G4a���5`N�"���B��y�r�aC捞X	���dJ�
O �'�f�5��͡m���*�툅)IL\��6Mx|���C!-��x�O�p�4���B��9��A���r�0����y�Ht
Es(����#�"E���X����[y�����S.��[����&Vvh�ժ��	l��[�!��`�!�$��">vm�CLC${&��Q�Ѫ�ڜ�c֤:�$X�7�� �*@�<AR�I �x�a�!|@zg��i�<qDJW�BY��X�"і�̕�MQ�*� -��3�@y����I	}\�H�؍�Ш��K���$ޕ�T��!I�!��h����+.:5�6�{?�l���Ә}�C�	�T)ԙڰ�h�@Yp#��_����Z�+=�Z����ѱ��pP	�4o��u�ǤߛE�)S"O, "!���q�"#��W�T���B p�%'n�!30�S��?I *A�FR� �F,��dL��	0��V�<i��B)x�2P����-���8ӧNyR	_7W�L��	��� �`��n��(4
��4�C�I'
]����瘿0��w�ƞ\g�C�	�h���xB�Z:M:����X.v�C�	�@<	G�� �B\B����FC�I,)ej���k�}N$�O�z*C�	|�tC �Pܵ�WM�	��B�	K�i	��0��	PnR�9�B�ɲ%� 6i� <Ebiӣ*P�7e\B�	\Mr� �"�/L\���u�S8G�XB�I,n��jS&�h�����/�hC�ɮ(�d�bT�FRT�z�F�'Mf8C�)� ��z����,��LJ �	.C�53"OD�s�<?�\(�����mD�E�"O��_-#5|��9�q "O,�AƁR�!h�ъ���j#p��"O�:� ?N\>�!R�;{�"O���	]��t�s��A���"Ox�K`��E�4)b#��0B����"Or5��A�9�L�S,�/	ĵ�"O�Q�QnAv���F��E�xH�U"OX���,W�J����@��4�( '"OVqK�<>�4{R�¸0ҍ�@"O �92�s�|��Q�s(�t�"O�<ah^&.]�T�ͤ;&~,��"OL��#NҨ�Х��Q{<8��"O�� �	(�`-���V�-���H1"O��4�;���a�18��!(�"O�aꂹ*ipwmE������m�s�<��D;@l"U�p�Bq��MWj�<�a.(X���4�t��Sí�\�<y�JU!g��CSL A��A��AZ�<颪J%{���= 8ڀ��U�<��g]u��9g���G��<C��P�<��e�0[��`lC�?�t�R�͔N�<IV#МJc�U��Ό(,�(xu*F�<���#5�M���\�k�:��-|�<A�B��3���*���))�ƨ���D�<�Q�S}0�Mr� ���zF$�F�<�J�#:�HY�$� �3�+T��2`	�p�l�2Á�bw&����?D��0��P�`9�PQ��#] $=D��؁ ��u�rx��)�&b����=D�$�&�ĸ*(���`O
(�lk�F$D���f�\�k����J8��I�U�6D�p�c�s�Ψ���կX;�9�8D����L�DN���/�^fj4D�(͒-{��42���$��ys2D��ҕ商n�42��:��G�2D�L�VD�;%pɹd�Ѳ[����2D���+͘/�Ψ��@Q8��7�0D��rfn�?�*���)�!?T�"e*D�y�ˡ6Ox��_VB�!E/?D�X1�M�pZ`�uX�8�` D��bF�=	l�� ��Y0$|	#!D��@��ͬi�)�cA9�� K3D�8n'���艱+G9,	�lcEO*D����Ӫ:���@�Ѽ]����%?D�谰�Qአo����y���?D����O�&]�g&��.�����=D�l;D�¬K�B ��$T.u�9ic�)D� �W$|C�
2��,��=��%D��$�.W
�@�EG���Fi�?���K�:T`�I>E��H.H���eM9y(�!S��� �!�ĔP�X��ڨ,s� �o3y���W�Lq�3�	y��y�k��U�����3y���F�ۙ�p>����m`��b�I��J!�c~���t��Y�����'��1K1k�$$����!���^ÄT���H�Y���+�&'��c?���^�T&�MXR�E�[�Dm��b#D���`�%M��ca�0v�z&�� H(8�:��s/O?������B�R<@�<��
�!�$U,	���#��4Z �d�&�"Si��Н:d�8լQ��'*�7(������rW4�P2��b8�T�`Ȼh�L�Y�'\�BL"G�/q^�:��.~�Dy���ԑ)Q&X���� �'�HpGy"�6���y�&ٜ�����@�2�؈Y%@��V4X��"O� ����� Ұ����ڽ=$$���k��d9R�*\
�ٗ���B�
�F����S�r���������y���66r���2<x���g����;���s�h����<�P��� �����[lI{��gx�Lk���'
�ca��d�R��oP�V>*��4)�ݟl[k�*
���	!Z��Q���2&:: �#� 4����d�s�I(�Ґ�?Q��Ү"��S�T�,���+$�v�<agE1y`�+�L�!M�`��ɖTܓW�����ʊ;-��Ë�iZ�#��݈���9b�4�8��J�c�s�a*Q���S��k$Ё�!˯A�hcf��0`F��B�
Ƞ�:P��9e�<��
�9��9��42 ��m�nr��'i`�i훍��Ϙ'�.2w��NY<X�B��/&!Z��@��p��TE'+qj���)��͠�Ʉ\���K�G�N@d���� �i�B��5,+�u�v�����,GĈ�4��!s�ɍ4�2@1i�	>�^�GBL<"=�� D�{%�S�6}̽��-^�l��i7��2\ߔ㞼3�"�i�J��N�u�O��a��a�&����"͒�|��#(O��Vc�7M.��3p� �̔�֠ǁv+�m��^=�{n�@;p�A��2ʓ ,�|�'��=x�IݢBo���SOÌ-�� �����d�9�8@�"#���JƦ�`r�����@�6>����Ұj$���D07�Q� c3��?�
�+��ӳ_�Y���
�y��ѕd�($��&Z�T�F~B@͚-��0�a��2�˖63]t��	
-}�D1#�O7�I)P���%h�.Z��T��b�&-���͟�y�����͚t� �]�F����d_�Zxx�f?�0f0Id�^0	_�iY�� 56��]�p��G�����\v[ LSCi�d�O��I�!E��TCF�K�.�T*:&a01�ȓ�΅��@��N+Ľ9ztk��h�N�"���
"W�͋s 64����6�	%`���{*[3���
@1�"<! b�K�P���G�A;�D�
�|j��Ǩ���D����B#~�@�����8��?�!$��UlL��%1hT����F�Lp���t?�C��.�p2$�+��O�.�NFN�1BE��6( T`.9|!�2�^�H���oq���q�\�E�ޠI��Db����6�j��p����LS��٧m&�O2�r�Ɲ6=�p'k�/2�"����'�l��چsR�l���^� ]b�J!J�(���
�0᮸����'��<�J�ް=AӁҭYt^}H��E�~S$H��MUL�W�D3Ճ̅I�b牎��Q�P
7V4�p�;L�d9+Q��f�P�T�V����'�t��iN28̸!G�ԀL������,��8k��Ol��L֯D?v���tKw��vMZ�~����.)�a�F4D�P�F��;�� 9�%��I���Gc�%@n\����f_H��'��̓
}��Exr���hj��f���-��g��Ӱ=��cS�X�c4��O|  $֊N2\��!6��q�"O��C���Z6y����;-::����L���1����h���R�� Mi
- �'C�	ʴ�"OQq F�(GF����؉1�^��� �gNX�b�OL��ע_צYa ��?����X�0���0��E�d
�m��(BB,8���P5"O��x��'h��4�#A�FO�lhbh��bm���O�IH���&�����'i��<��Oh2$�ws�l�t��-SHd�1O��EP�'�f4Q�`�^�hs��8]g�$�$��u��0��K�T���e�Oub a��N�'� ęWf�5(}:9Ag%�87�*U��)y6�e�:4�>}���@�xvE`�3?��]�H�!H�$�Wsj��sN>�O܍�El.{��:�/��F�I��|�Q�J�yؓ�ܛ[Ȣ��'+@�F�
�(�D�ti��q)F �@@ӊaaLP���ϭ�y���(-���(a��V�����)ġ�"�]���eXQ�U�1|���=���&���wg
u�e��-l���G��x��	�'�����T(<]t �$�I�O��)��8�X����M���Ҵ�ޙg ����/Uk�'��\�k�O�hѢ�'u�)yϓN�d���%}�)T�̈́1>��e��}���K��N�ؠ��]�H@�w�>�ON��0�װ��Y��@6Md��0��|� [7Nc�� �-���v��ޔ	�}���H�&�&���B���w~a����y�ľ|�>t2e
�lCtp`@6JyJ��7H�Q�$��&G�� `����� a�Eλqx�G�נ:a��R�ڵE���<� :��?�$9;��_��M�^��`$K��]�����ʉ�e�"UC�G��H"�R�8/|;p#Ѩ3���#-O� p�A�A�����O�Q�s�ٳgDX���$&n�eK��=�)[f�%�O��⃊>z����w�H��>�s��%��-�k��= Dt@�現?%nlz�.=jL�`>9�F�'4����V�<� �x��_��~�	s��)k�ᘡnI������LG�2����`��q�JM3���y�/J#82FCR.�r$ h��Px2�G�z���S�O�"D�T�,O<ƙr�V9=*:��肵L�"Ԣ�*B�b�G|2�T|�h�� `eؙ���E4�p<)bU�+��Q7*V��eb��;�M���;K�T��ω0K������X6*�,���_�e� xjB�8�T���D�\��Zs
�8'�	u���3�IG&��Շ�sPT�'Y!pA�$D�;ٶ��v(ʹ
��Ɇ�x���`$&d✌`%�N�����g�bGFP:�	R���k�Xh�;�J$
6:O�x�A�ӌq<h���_�D���&O�x	t�Ѹ�����G�)��[$	�C��+�Oѝh7f�1b[<F��q$1�A�����̭`��
1`�C�`1nXd���ĉ7)Vh����dάA���K�6X`�� �+��2d�L(����-�E�'�6LH�A@*)�쬦O�(Xpo �8�I�G��?_4������,�j�	`�Ax����=^���<�.�8Fd��R"܇.�|�r$X�t�UG�s��¥��`>Q�#͜�.�(�X��C�y#$5�q�=��Y��+�g*:�͓�ң|�',�%�G�E�wx9Pi�ts(8�FZ��@�^k���@�:��D��d����ݾ<��(Z�-�n�YF��*����C��4�џ�: $2,<P�S�O�0�&�1�۹���D;0���F~"��k�Ľ`�O \�e e���c3�\�p{`{���3���3o�w����O��qР�J�@��`Cʑ�3
|�1�b/0�9G���ŒWĵiu P.�P�Jd/��䕀C[�X"��?om���0�Y*��̆B H�A`_��!��G"�HJ�G9�`�һ=n$��A�"�򤂸I���1�/��$��A)Č�FDF�p�ƭ8o]CB�2dܧB.(yʒE�3�8!zt�W�z�q��mR&/^HL �'�*��� �5ɈE�L�yu\l	Ó���`���:b��'˜ii�͖E�JP�թ�0@��T��'�$TtK��gi5Q�	ͿmU�O�,z�
��~ٮ�'��?��ώiVH�ae!7ql-lRS�<1r�S8~��j5�D".߶5���W�<�� 7Ez�ȱƣN�3C�5)G�R�<�'�M'e�0ɡ�K���0�E�<�)�aJ|�H��C/��� k�<Q�� Rrb ��oXH�Hy��b�<��ŗ�4|"�҄��`�M���PQ�<��CF�tц�� ¢�B@Q�<�eG��T��H4X)�`i��i�<I����S@hpzqˆ�5x�s�FN�<���C8V�rD���.p����S�<�rl��w��]�4ʜ M�����U�<1p�P*Kb�1������A$S�<���R�1j=��*^0$�$t(���L�<y�O�w� �d ��L'n�2���s�<�wU�w�bf�Z�A��Y��Jq�<)�i�>G��`A	0W,j���Bn�<Q2����$kV�Ѷ�l���d�<I6%Qm�F�BO�?nY[� Ic�<i׫�8s~��,��=
9ˑ��X�<iA�ÐZ����M_���,���AV�<��!�}3�D��.��k"B ���	L�<a�eJ-M�5��MY�$'�A�c(MT�<YӁ�B�R��0ϒ�x ��;dR�<�R�[�䝀�%1�M���SI�<y'��c!���&�^9a����F�<�� �3&�Z<�G�Lb�Z≚E�<!G��Tת����g“�m�C�<�Պ�4_��L0�^�X��ЪE�<Q��[�A~��I��] ��;���h�<� N�d`f�A'�_�ij�	���d�<��G.#<"%�g����9�w�x�<�BO;A��Atd��a����A�z�<	�bQ�v�����eL~�z�,Bi�<���0a����F��P:Ĳ�a�k�<�t���|�䆓TE�̪���J�<�  �s3��T�dH��c[�1����"O�`"ࡐ�t(��1g��c�^d�&"O$�еg�5gڔ�I��\U�z�Xp"O�l�U�O�:��[�٧S{�*@"OBe`%�tr<��E��e��"Of<1��jI|ܙ�n��p&�F"Ofd;P�7Oqh�P�:H�e"O9W�P�p�K�)L���#"Oh8	���S��(�LBȆ# "O�Xx�fX�} ���
�l�$R�"O�!z�N�+���� �X3y���0U"O ��g	�TF�=����E��9z"O�%&JrT��S˖�7Vr��C"On�b$
�]��lqP�B!6��%�#"O��!@�:� ���ΔSm�}C�"O`tѡ�G	Y��hso\>K��I&"OFs���?b`(HΗQ1�5D�l�A�O����&��>e�6p��$D����Mp�a'�!L2(�*O.�!�F�$(�Y�Eb�\q` K"O�e�0�R4-Y��Z�B?mL�W"OT��C��J��4�ʥa��*c"O�kt@]���t �!E�e⭚7"O��i#	θ(��)�2-��iX
A��"O����쁁��)gL� @�=A6"O
 %�A{8�'+֡}�����"Omb� �'PP}��%�7)&���"O(���Gǥu����D=%�I�"O�ِ��K�2슀I%���"O ���� vޥ��C�6T���"O�q�B���tZ����l%jCeq�"O��y"�ɤ\x��p�@�K��t"O�aꠤ��a&8 b!�)�"�"O�����|�������$LH��7G@<�Űw)
+O�\H�>E���/iH��F%ڑo��D��H�y���:hU��L�)�'@V��B��ќ�ܹ�Rl@~1�pΓ�?���ݛ-�6���O�˧n_6��/�Ũ��w�	�����@�pl�A��}֜��S�s��O9�Xa�@�)9���PZ�F��ѻ��x�Q���<�}�E�4*���zbgH9Ek2aҷ��[y�[�`�<E�ԧ[u*nbr���u��k$o��?Y�O�c��'�� nl�i���ڸA�th۰�ېW��X�q�<١M�>� ÒC>	�O�,�$�:���嬴�v�O� �''��
ӓ-�xVl�1th���=�n-�g�1Ol��%&�)@���"N̪e!��ճ#�B�ӓ"Q:/�!C4���'!�$	�+j���.��+� 	* "��%	!���)���J��'Ƙ�:堔�*�!���}�`���n�\`����"	�k�!�F7=��K$J	
cBT!��U!9rh���S>a�B0�P����Ț{/�"��j��	�'�f�ź��T>Qc_>5���_���"��B��"�
^�L�,��D1D���
_w�$!��S��t�9�'��zE���y���A�'z�����z�՘��^>�CS.D�s�.��&g�@��b�G�4�@ 27�B/;�*mzF*�+'z��)� s��Y���&�BL���M�/8����_�4]�B�<m�x��O{�>U��CU��{ABϩ	��r��E�?�dX� �8%���`)_�<E�DfV�v��|���b�<b&E�7	ed1b�O���'��M��ӯW��� ���>'�Z��Fb��HOL�2a���Ҹ��OS��b�D~��ye�ڋ]�P�i�O��kD�K���=�ǨB�j@,(�|��1ӥ�}�<Q�ɏxh�d�ŗBz��J�z�<�8���`���d�$�B �J�<Q�P0��T��@��A�h��3�RF�<��69�R�H%kSj�avfX~�<�bJ�#�R���cʹ"m���F'�~�<� ̙y��O?IDR�ȧ�i(dX�"O��঩бU��� i7	����"O8�1 J�?�j��Wɞ�{�й�"OP�5�ŤA���BQ�Х$�8)�"O��I����*�W�Ůb��LKc�PM�<����YP�K0j�*X�(��N�H�<��A2O�Ѐ�2e�R�8��X�<ID�ԎO0� � C�&����W�<�)�?���ta��������Z�<Q�g�%5�h�h0�[���q��&QB�<	��O/b�� � ��,)�L�0�{�<�Roȓ ����OD(<�vqT!�p�<�V��s�ZaC�&W:?qȸ{R R�<e�5'��s�	�3"�X�S�dMT�<��d�'*�Aۡj��p�hH[�Xi�<�Tn�
��5��i��xF��%�Hc�<y4�I�^X����E4�({�o_e�<���G�#��j����}��(h�^�<I�GK'{�<p�M�� ����Ň�O�<a"ȓf��k���@��Ta��O�<ٵJ�T�,)�1$��,l��iAI�<�݈w�LJ�H�h�
TG,�i�<I���"n�Yס>~B��$�a�<)�DD;O�@��k
7g��(yAe�`�<�R��K.����+9��e�D�x�<�� ��9
P�ԤB�{��#��u�<�$kX�*J0$�����sh���l�l�<�AI��<.�%���>�d�@eQ�<�я��Y���+w�Γz����ly�<I���#�~�bPB��v9��ot�<��j%W�>	 rb�G��:W� x�<����}���q�@�r��^{�<9��?B�<9�����TL���¨�s�<��U�[�r"�!A�p\����&Dn�<�F)YYC�@��
S-wY����t�<qb� �N@���@�A�
 �ѣBx�<��D�2x��um��No�ai��k�<��J�4K���� -��w�
��Ѫ[�<	���^?`)9T#�"S�H����Y�<Y��فb��t���Mfr�IE�}�<IG� �U��͒���?@��x�P�P{�<��N��%l�۰D?q��x�c͝p�<���GX<��G�f����@Ut�<��jP�����ŅTP,�@�p�<�TΉPC�FR6?a��b��Zf�<��c�r��89��׭
��	Vb�<���UL%p��ݩo��A�f�V�<Y���)$��IG�M$P�x��	V�<�Sm�-a`jŊD\�\JirCM�P�<U&�<(l�@�&)H���  ��M�<��j��֣O�o@@�iT'	^�<	R ��~�� r2W6I�b���̚\�<A�c�,{R�׽^(�I�n�@�<A���RL�8��!V J��C䉁���o0���J4�
zF�C�I67�J�ZsNF�Z�����8�0C��#[{6زGF�@�y��̒�vq�B䉴�^� 7�δaO�abVE�5k�B�I6֊�1��~���u��?��C䉍a���Gx�%��D.,��C�I 
9b�Js�M�Ą��q��*0%�C�ɢj��'��V�V���M�Y(fC�ɡy�8�(@�]�B�,��g�
}�B�{t �a�>"�I�`Ά�v<B�)� �I��NA�D�Lt���(2|�K�"O|$W�^������#M(*�Ũ�"O����j������-�D9HQ"O�c���+Nȱ�L�==��9T"Oh�p���/r׺�c�F�=�͈v"O�m�aE(|�p5eE�XX�i��"O>a�EaP�"�D�l����d"O,$zb"G��Љ�m��JØ��3"OpK�`]�2~���6�5[�,��"O�E/�^/LQ0�'���`�"O��F�ܪ5iT1y�H�V(&Л�"O����3=`
Y�e�f�:��f"O|�t�X�ۮ4ڱ��0��eyq"O���ŉ��k���IՄ�$(��=�E"OXy.��\q��B�	J�bz�4�#"O�����k��j��[pP)�"OH�C�4I|@�6o��X��	�"O8���I��PH8�'����(d"O&�з�F�H,�(�(��q��ٹ�"O2}�񋊔c:T���(�~��5�"O2�*�ߕNʶɵ�O���q�"O�x: �YJ!��0�)]^��Xۄ"ON	!���1M��(j@2\�h�K�"O�}@wN��E��ʔ�L�[�9�"O��Ks�ȗ"��+�J�r��|
�"O\��b�c��27mB&^K2$`�"O�tbT�g�0QǫÚ_H�3"O4�@�N$Dh�� �
W���"O�0�J�Sf��c��^�铷"O^a���EcD��@	R�f*�4"O�;R�G c],8���O��� ��"O��1 'I�}�lm�aAML����"O=80��+Ш�r��R
B
P`�"O���`MM'Q�
�#�n��b,&L �"OH��Q3YyTuS��_6\)�X��"O<mX�)�:,c��{� [X��t��"Ob}+உ�1�~0 @�R���J "O����MT�ǐ�QE�Q���̉�"O�U����-EY^I-ѭt*$H�"OJ�#��8+:}�0n!y&�D�Q"O���#�6m�8���ؿR�0��"Ozݡ��ZzDH �C�k�v��"O���ГC�����B=+T�\��"OZ�*&�Ɇt�d��a�9>M�t"O\���/�92-4�q`��2[D���"O���1��~=@)O_�vT���6"O` c�ְQ���sÆkN(�6"Op��"��V{^����/c
P�"Ol��'�;d�{�ia�*"On��.Wx}P�[s��z�����"O�-��DŘ~��`�T��2�� �@"O���K�1^l��
�{�<�H�"Oڰ�5Ɨ52*��@炖cbx��5"O�U�pD6k��]!��DPa�"O�y��gҥ,�F�O�az#�"O��)�$�"�y�R5[]Z�A&"O���z�z�H��$l|Hh�"O�Y@獟�r�B Cd͙�#O�:"O�t��D��R�)S�+��C��# "O̝@!� A��l���̜!�"ODQp�ъ���Ѭ��I�8I�5"O�ѵ��|�T	��W�l���'*O-�C�,{�=I"��hW
���'{��&��t�"��P�p�J��� �A�d6R_$�b��5g>�x�R"O�=�k<byBF�O> �"Ont r��iφ*�%�t ��Q"O�����#P�\p���i�hC�"O4Y����@ꦇ�_�|��3�Gl�<a�m�5Z\m�v�ʳM
��PA@�<q@LT4M��������=tu4"�~�<g�	U�z�Cҟ(T@TC�{�<Icd��_���@K�C�z]`vd�c�<I�j�V�x���H׼9����È�_�<�%��KO쑢fZ�M:V谑nLT�<y�� ) �xq္�$�
�P�<��Dpz�ذ�X!�gaTO�<�D	a�`]��˭]��(�@�E�<Y[�� �w��/q�I��	�P4
B�I�n�Z��u�P�r�	#�� ��C�I�9�h�c�������3$_�C�	7f)�E�wf�H���{���,�ZC�	�1�P1$@&Z�U�׎B�]�$C䉐?@��aD�	��I1B+��T>C�I�v���H��2]��h6ˊ�6C�I�
�6���8c��!��#���B�.I��4�U�XQJ�(֧�4"r�B�	��}���~f��c�Bb�B�	�)����@ZcF���FZ��B��7���s����=i�a���B	O��C䉃B
�Q�js������C�	���t�p'
�7�����p�C��=S".����I�y�`bW(�^C�I-���p����$�T�vN�B�I�}r�Dra���/�l]��Q":�zB�Ʉ/<x�S啧/��ãN��B䉉2N�r�^?P�~�`狇�:IB䉑/^�B��[�\x��cf�C䉬W�^�c#aU�)�8�3>_��C��0=x ��GÎ5
�i���1ȗ"O�Pr��Ryv��ҕM	�1�DZ�"O�$#f�͇E�+��3g.t٤"OT�#����*�Ȁ�6�L��"O�=z%LϿ{����D�ęP)�"O4mKӡ�/�p09�ė�8�N!��"O�� �+[G������iX�"Oh�� +�F��[�����`�"Op��Eo��^fl|K�^�y�JI�"O�(��;k�����Cm�}��"O��`��S�ʹ���*TW<0�"O�Q�q�A93�@y�"��e��a2�"OƈH��8 掌��%��b�Ry�"O�a�*@�[jT"����}j�"O�� �&�#)�(�H��M�J8�4�f"O&��HĹJ��m�ǆ�!>H3w"O��cn5Z�AhR@��GZ���"O&�y	�LP���I�/	��j�"O��`M�L�P �]6gҾI�"O�	�l�������: �i�"O�Q���r�����  �"A"ON�;LP\� �[F���j�08"O2l��j�`Ԡ��ǘ�@�k�"O��	&�ѻ�)�'�<��"Oh��6LF�Z�2�{�蔶<���"O�\9Gn�A q�C,S��A�"O�Q��c,8'����^�}|�hQ"O�����a
��Zo�1�"ON���   ��   W  I  �  _!  %*  �4  @  �K  �V  =b  �j  xu  �~  �  �  !�  ��  ͨ  �  S�  ��  ��  9�  {�  ��   �  B�  ��  ��  
�  N�  �  �  X � �  �' �- 5 �; �B #N �U �\ g �n %v g| �� t� �  `� u�	����Zv	C�'ln\�0�Oz+��D��`�2T(���OĴ�^��?Y�+��?�����,+l5X�	�[®��d&N�Y�P�����F��t�T
%�iR���oh�I�%F��)�Z���I����Ud=~2h0���R)��k� !���ÁC�u�h`D�P�wb�ح;^�,0���H������ud�1p�<� �Ҽ.j"� �&�I�0���u��0U�ͷ-��un��n����ݟ8�����	&;֜�p�K��.w (��b�z�����(DZ��I��M�.OD��P
���'"�;�ꀫ�>,B�H����0k��'PR�'x�]��w�t�M�'�?	��4M^.�ä���t�������HOR�F{�i�4#�X�\�M9���\[���"�>�����.,
���O�=�c̧)�fAXaA�%��@w�')"�''�'Z�	�ܔOU��ًq�!pa�b�|8肤K��bG�O�6�ɦ!Cڴ�?���i�\6- ͦ��ٴS�J�۴�_Z�.mN�i�pb�'/��I�O��$ <l�8�d��S���O���Y���~�4�x!��X��!jמ�����k�`���#��6N���	�?���6��KdFx���I_�ѧ��3�MCu�C
w����&	�:�ڑ0�|�,�-�_w&7������4X�z� DbA�AUpID�]�_�и��	�����X��o�8�M{��i0H��q��,艋��G]0���[n��1hU�+�	U�J1"�bY�e#�+V尢�q��\m:�M�E�]��t��h��nV8A�i�m��Y�R�晱�hV�q��榽�f �3um���õN��}�I�ٟ��?�3���M���:D�ҼZ\@�(����?وb�'{�[d��6MCt������fĪ�tDO�6C� s�D�}�����O�l��O���b>�w�iO0��/��	�CT��ұ�Ƅ. `41���"z����ܖ�M���
Cd:���O��
�J
*I��R�ϰk����P�'VTI:��?�O6�q'*H�ڮ!��tP���'��	J���O�`i�&�H>W'�;b��. p$Q��
k��k�B��������*��?1�I�����]��$E�Z�V ȇ:��B�z\���훚O5.���bŊ{��B��$7�v��1o��$.P8e�B���%c|�Y�U�dsC�� I�> ɦi�/x��� `MA�C�ɳ{����-�l�u� K=|=�4oZ�X�I�d��9�
1�	����Iҟ�� =�v,X�&]�.�ɻc��x;��p��ɟ!k i�� S&%!&��F�C�D�O�J<%�|�5LF=SH^�WoZ&����ìϲe��t2��I@�NQ@R

�<�Z|R�jKa�t�1�"��w���Q�C�:V�	�C�֤���i��˓J+�4���?�����@�dg��_�Ra��Q�:�V�J>����?I*O~p�O��Pi�O_T�2��1
r,�8�Q5"�p��?Y�X���'C�韄�O��\ZD�T�ual���hE�w�XL�)O(xJ��'��B�֠u��ZT���3�ax	�'$�Őզ2t��r��#�Z���'�ڸ��Ȅ`�p�L��VH�	�'����ȋ,�tC��i|�;�'g`|j��� ER�"P��"<w���
�h� �+��?�c{b|���o~��r@I�4�s��?�e�@(�?!���?	�c\�n�L8+CKK��V�J�w\��r���+d�@�S`��=&�D�	Ó]	��b4O�H���%�ϑ ����kZZn�
�n̻?Eh|X�	����Ol���'��6�����I*���nT�lyaw�*PP0x�I��	ԟ���a�SR̓SR����,���B�+`� ���'��}rk�X�QoRwC�T!���	y+@��NŦ�<Y�4�)����O��t��HD�%%2�s��D��tA�'"O<�ԥ���x����~��"O��⛆#A��Z���n�!p�"O�Q��b�k���q�<<� �i"Oʐ;���:ph �#��}R6"O�Hqec;"�8��/D9*H�ՍhӢ��O����&a1B�Ol���O.�����9# �:'P��1!�c�4��b�S�#J�(�#������
ОjP,ėO��⟨��� fS�Aqs�N�O��Ap�H��,>���r�x����c>c���ժ6�L�iPI�a����O��'���`���b�'��4���/O�eI� ǼEP���ې!�$ۑG��D��@֑>I� ���2�	��Mˤ�i)ɧ���O剫C%����'=�h}�r�ǝu2H� 2�� ]��y�	��d��͟��\w�"�'9�i �H����g��r�f`!���2c>�xkpO8�$a�0T��z���Y� @p�c�!���0P���D�6Ȅ���D�H%��b��'L���ĝ�S���V�E?�*b�5T�!�$�`��ɛ��B�.���"/�w��'L7m>����h7��O�B��-Al��8Qg����1�I�'RC��'��|`��'�22�`	��.F�Iq�nѼfM�6�#� dɢ�<-=�p���-������:�<�\P	!+�;�& �फ़�MP�N�|��a���<J�Ked#0�}�
ڲ ��O^M[�'K���T�ǭҖfW"�9F+̢~tp���E?�D,�O��u��LIt���yE8���'%�d_��8�#��,>d�СrB���Z�lr�'Hȟ0������O��uZ��'����T��I���)�	h$ac��'u�*�h8F���>5�j��cZ��NA����i�qE�x d��#�������	�Y3~Y�`���Wm޽�4���?���]w$LB4W>��a�^���7i��V%N=���-M��'�>ΓO���2��*JF�4(>��VB4D�<R����B������p�>�?���S4c��m�!��K;"<��/��W����O��dk�������~���$�O��$�O��]�gP�RVJF�f�L<R��3x��3S̸xmZ]EU��g�Ţ��x!���#��7۸5�p!�:@j�u��E���A�4?-��IM�`��OH��� >�yG�A]��y��ܷ}�@$�;�?A�O*0�0�'���.q8l32f��N:�5�`Ğ�G��0�ȓ]~�:B��t~@�kT!fn��ЭO"]Dz�OE�Y�x�RI�&B���3F鞆2�)Q�b�4j������	ğ��I�����O��$��Kn��Q�E���M� �#��u�P
-
�T;��U?m����*���	��QP�� F̴aGٽ:-�,���P�&��,,��<a�f��2e�|����c�f�i�Lk��I� ޴�?�+OZ��;�I�LK�s� �2�ᒋ�#t�$��z<����{���[pΏ/[6�s�XU�ɗ�M{�i$剫F�� s�O(�d�&�T��wU�FtS�J�q�\�D�O���L�O���i>��4�\�>��R�	G�@`lZ�]�J�à�I� �(%��j�*�؉��I�\8�e�N�=h�*�,w�
M3�nN7w�"U0�D�������-C���O�Y�W��	�	����'���#S���c�))CW�0�L>1����CE��*Jݺ�]�ua�a���	�?�g��W���d�3;������ �'g�����'��'���2pE:�	�W.�(�BLZ<ґ�Ћ�9�����@�'��*�H�CLӫ`O���S��?ep�.Bs�� ��L��Bl�R�7?�ĂAq�9�׷;o��1���,+�pP��.�^����J!<����\,��OZ�}ʜ'�L�J�N��?D��ʤ�%}��,)�'��)�C�G-]�%k��/wb�9[��D�^�Oc����!�9pL��
҉GGJ��"�i>��'���T�cO&0�7�'���'�25�QE��p$�k�g����8eH`6�;Z�0	"�ӍN�`�1�1O�L*q�A���P��o�>y��%`+�>"eԀ�	Î\��Q�Dl��2�1�1O�qo�
"�ӕ��  �H$�y�ٔ'*�q����'��'ex,"�Ma�����!�g�Q��"O4 ��Y�9�pQZ�b��GUڐh�U��9���馽�	N~����)��t�#ˋ�m��c��<��P�P�|�Ӽm���� V��Ea�� �yr��?#-]���Y���K���y�HV�9��uX� �9�T�J�y���|-��h��Y�C��1���yB�h���y�,��7x�1B����>ɵ�p?�a`A�B|`� ��N!�U��K�<i�j����C�i-�)"�$*�y���90c�m�"�̨2�z�W����yB�ؕm߈ Gi��}�f��׭�=�y���I�8���\>p�P]@��^*�y�ԲL6(U����,b!�"O��hO x�B�Ӛ]a�re
�2lY�4�ӏ�V0�C�Ʉ/CL�#Es��,���:3:�C�ɂb��8��ONI�t�w�í9��C�I�G�@d80l׺yfr0����+N̆C�t.hEO�Kb�
1JR��ZC�ɟ.`.|��M ��8(�&���|���$$�"~�P!��<�&,w�$��b� �=�y"	G=py+�x�b1�y��vXx��O����yB�,<,��e
§zkj�3�߾�yBY:�	W�:b{
�*$D��y�nA����5��T�Z�pS�[ ��d	7��|R,֔t&�`*�+�E�l�y�!B��y
� �<��T�9R�!�(U�Y�$Q�"O��B�o�7|v�pE�o� b�"Ox�&�8<G*9��+}0�$"O`0�PJ�W�j�3R$ɣ/h �)u�'��@��'���+����M�����%�����'�*U��ӳ�&�l���*�
�'������K���5Oߓ
&x��'.�  p՜+���X%�
9mƞ�a�'���f�T._"�D�T���V���'��<��'��CjD�P�iL������I�E�Q?Ź��V����
�(� q�`�q:D�P1�&ď;(����E�Q\� S��5D���դY��ɤ�:X�ѕM3D�,QH��N� ��?a�F�o�j�<i��ȈC����i����#HTC�ɫo��U@�-Q�N ���0�x�`�d��K#�"~��o��c���J5�?4�3�M/�y�*ëcv�T�!{�&xcsG�,�y��0"Κh8�&%B�h�k�m)�yB^< *�H��#%�����
�yF\�wfV�F.Ҟs2|i���y�P#$�,����lx�E�1JE���%D��|�� 7δ�"iN
`;2��g6�y�i�,�� ��X�i�\��m�	�y��� R6�1�߾*����h��y���F��E9f�Ȧ(,^h#�O���y��֙@D�!�ě!����a����>Q�l?QAʎ�!�Tᠤ*��((h(��Oi�<��a�{b~l+�o�j�-���g�<�vK�E�,��G���LD)!��w�<���P�n���ē$�*�P	K�<�t3b�QP�`��7G�F�<�U�ރ6��E��@Y�Dw��K�!Dj�'V��C��I'D�d�`i@c�FY��CD$]A��Da�I��ተzX�P"�׬�yb�O�%�\,x�(�yjTh�2�Q��y��L��]�"��s�^(��˫�y��X�=씕tnֹ�t�B�L[��y�LS^D$�"�����|J�IV��?��MP����x��6:7������L�0���!D�P�uiW?>���'E�&���c%%>D�|!po&%���e��%��6EP{�<��;t�bqi�+�OD���UO�<�t*��)�,k�n�"�4=���e�<I�Ř+^�>�KFa߶m�$
��dyr��:�p>)�Cͬ/?L��%��[�$�IqcSI�<��?y�tɧ��<�5�橅I�<At�� s�%��+�_ƈE��M�<Y�J�|�%��#�3i�����~�<)����2�	5b��iYu/�xx�������H����*2Z�	a*S�e�h�J:D����k�Y��}�7�ϝ@�*<�$�9D�(тQ�kt�q1G�#[n0��E�4D��a���Br��F(3�	�!1D�L(��r���2�_K����`�.D�$�5D���%�ܫJ�����-�H���F�T%څNnj�`$ 
1Z	��v��	�y���)�]R`�{�⤙ŠF��yM܇7cphj�EW?m$\����y↑t��C�o�%cR�\��̄��y���u�N���h���#em.�y�H�vQ��h��S��lU�Z�?��*�r���������C9;��G�S�"��S..D�L+S��w��d�>�J��-D�� ��9���?'���_}a"O�xȣa�1n���aF�3F��"O�["[�4�� �A�/1~���"OH�A��-S~���!�=CsT��6E �O���dG� ��YJ�K=w=BD0�"O�����/ ����i�*�8%��"O�0�R��͚�g�1�y�'�.D��S��ڗ�HP�!��{�r�)�d,D��!񈝤K��H���U�nY��&�O��`�O8Hx5�F�a��%z	9YA���`"O�	�m�xp�h�M���8bB"O��W�'�V=bጁ�<�83�"O��0���"��#3���["O����c͒H�^D�%�/���x�"O�eH��ާ*NbM��嚑i.91��	�	��~Rf�>o2\ɥN��b�<0YD��U�<�V��2S�����+��̰�P�<��/�0�T�;�Y(4�ԉ���J�<�'A�-�hj��&�
4���W`�<Y�HP&�I��Ιyy2�҇�r�<aD��
{펍�cBܔ F`:����PK '�S�O+
�	!l�Y�Niq��e�!�"OBI����W�� �`_��@Q�"O�X�����3v!Y@�L+?κ�X@"ON�YCfְ/̊�q����u�B\��"OF��ХJ2ZLp ��8��5�@"Of���	3sb�𱳈�2Cq��#Y�t�4(1�ORY���5N~>d��J��e��"O4�w火B�	zХC0�.���'�Rh�0��6��Q2�N�.r"N�A�'zȉs�\y,��3O 9et�9�'� ��#��*	��D{C'S�y03�����
���@Ԉ�"x�6�郍�9
��<��;�D1��`
��7Z�'�<��s�vu�%��3;F�p�7�=k]V���)sY��*/3�ZE���Gb��ȓ���!+�x\�i��Ӹ�脆�A;L,��/� ��l)�n��SHr�G{���쨟�����c^]8�Mښ �	��"OV0	��O/�]ò�=ϰabB"O��k�F�n��c��%)�����"O�p�����A�6���@��;�"O�i�@ �"|Q��CCi�'Z"�eJ�"O��i!��-h^�Yi��F������'�F y���/�*��OZL}�T�!ix>��ȓN�̘�W�T�"��d!�$[����.�e2c�4 wd��6oE H����PƢ]�2���jV�rӈ�|5��ȓ"Q��(�(�-9��e2V��j�nu�ȓ���A���	4��c���zB<��'�.��	�D =a�1Sf��ԊUU��x�ȓ,����J�	�n-xbH�4QH|���/�b�ABf�^��pʇ�~��}��A�f�A�V��t�s�F��p�ȓG:�xb��"5��0C�,A�v����	�V�I�pV� fbU��vq����/ĪB�	�oӂb� /,��@ ��B�	��<�L�.A�D����F7�B��!i���H� ��I�ֽ���K1? .C� 1�"� %R+gh�հG懎O�C�I'?�Lрj
�Y'��;T��'��=�%&P^�O��$��-E�A��я�|�3�'LF̒2�]*/u*�(�#�Rx���
�'��+��^�YJ��çeMR�N�q	��� <IG�Z�t�B͚G�Q���""O\D�%�'�⭹V�;�8��"O��!5!߹}B�p�\� iX��'�` ����S*��qϏ#j������[�j��Ԇ�k�h|�f��*7+ư�!�H�K���ȓC*Qhf�F�!���U	�)j�\��W��C��W�,�$m�/�:*�����%~p���� �*��}��8)J%8�\1�@�P�n�8�':���d����I	c<�a�Ā�i�<��ȓM
�l��D�;v���v�ںK�i�ȓi�x�G��7�2p�L:>��%�ȓv�F]97艆{�8P��4M> U��L%��Cu,�1Pԛb`��l^���I8��ɷAF���Z\ǺE B�AAC�I#`ÐTK!�_��ݲ���z�C�	�T�v�I��4`��P��2� C�IJ�4�%-�N��t,��jd�B�I�c��$�"TΌ���_�	�<B�ɷmU��Y� �GJ5ڷ���H�=���j�O�ҁ�%YS���Y�Q�-���'��Zs�?PD�X�&�Y�7<ł�'�:Y�	���h%f0$��x�''4���i��s�^���ܝ���yRk(���8��
=�Q+'���y����&��|J�7����.���?��X������B��Оh*�d�O�����3L?D��i��0^<U�4��K�����>D�0ʆBEd���u`��S�XJ�#>D��#%�2<��p�U�:�����3�y�N�g��y��3#�2/����x���4PxikA#Z�x$� s�[$w"�>Q���K�󄋿x@ϓed����OV��A��//]F�9"�z	ThQ�!�OF� �E�O��D�OR��AYg~�8C��L)� �'u>%�Ƣ�a������ݺqTv6+(�l����j�el:􈎝2���S*t���j'��#���(��Ì#XF">q��OD�d)擆��Q_�� f�Z�f���S�|��	�'��9&�;��	���b����$eyr�ۂ7��	��>2@aC����D/s�����O
���|�ԥ^��?I�������X,Z(�b���*9:y���V%3d���
y��%�=/ܛև�~���4�K4.�]ʔ��:^!B�#U	�y2/�8xF�0����\�1�C�i/�9"��K�dH������P�E:�|�sT��p,���"0OP���'⑟��^�M��@s���BPb��RC\��!��O@�SBK��Աf����D{�l;�'xd��"�O9T3�|Pd��+��1���?Q�3� (��Ã�?a��?������^[B���*�<^>��&��6+Ӣ�I��ٷʛve�	��mЗ�V���C�xb�!�g�EY���.\h��@���MàO"0��a�$����铸}8����a�<!d� d�!�w㛄��@���ZR~�7�?��hO��	�1�ZT�
9�R�㑯Կ<��B�I+E�.4s�BёzP����?_)���L�����'��	=!�E,LL��&<Rg ���I	*D�3w�Dş��������?�	�,�'+.x�dŀ�;��q%`�.
�\�vh�e���)�anƉ�Aå[鑟h����x����s��ay����a�542�{� �,P x�e�{y��2ش�M���Ds?�u�"��x9��^�m?������hO�#>�B�h2�)�@�6��	i�<�@����d	�&�RJl9�sB�gyҧdӐ��<�4�±=%��ğ�Χ�P�+s��V�����ɟvH��	<���˟|�ɻ%����`�ŋe�hi5��'������X����WBŨ~9
q��ɁÂ����M�j��y֍99}��pXwfl���W%s���Sem��K�.�z1�i����'p��I $g�%	�W-z�Q`R�	5!*��o���ӥ؋ظ���V!)k�����(�O9�'4�p"DOE�8�T�Z.<8R)O�H!��O���O�ʧ6�R�h��?1F��by��k	F�p9X��ќ�?���{%�q�0!�6�BHI��?5�|�rge|��-� ~!d�*U��<�DGɪ>�°��^�dԋ�Aˆ��ݺ{�����\'�l*�(Rc��YA�ő�y���@��O~J~z�O� ��" Cx���3͝5'���9�"O��Æ��(V&%�v������s�	�ȟR�1˃.Ҏ����	19�tu)���Op���O����	�45���ON�D�Ov���O �맨�3���`U#o����S��"N����I�z���Ej�.��g�'خ�9�M�>L]1��
�z��(`�F�d��&وW�v�������	K��!�V%ڡJ~	�GE
1I��@2�`�	؟ E{�4OT=ȗ��:%66Y)�g^�EOLT��"Ot!C��@�`G	V;����'�b"=�'�?�(OD��4@țf�>Lb�-)Ȱ��w@҇SŲȑ��O��D�O����<���O���d��5ξ
&ȡ�1��2���@㐉riu�&*�ڥ#�͐;��O�(� N� ���R��>�41���Ĭ��Az��Y!v� �R�_�>��Po&���?��O˟(j!G�,XP)I2G�V��с$�ß G{��I�$2c���w��pI@��"�B�I!݊9�i�:��Q��FT��.��'+剑i�xy��4�?����d���wV��0EC��_$� ��?�G��?���?�g��?qMFC�;jJ p���EXZ�U*��V�p�`��O.�@MK�u�
���̛.
˧}��`����J�Y"�\��qD|�O]��?���Ɏ:ar4��I<_78��`��Z�!�'4&�ㆄ§w��8�	�\9�}b�<ق)�,{���p���L�)
s+My��'2�|ʟ��f��3�;}��4D�'u��$�ǌ��l��HV�߸'�ў�3�)��}@��Xd�Lc5,:��Ԧ�$��x����X�s���P���4�[��	�|�7�Oց���f���O�O����n��u�{f��9*�@�P/�9&���%�n8l����0礑����W�}��������E�c���%�*x�	���i����������<�^w9R�'��D�'M�$�5&��Yq�OO�SJ��R7�^/~�MkR�'���ګy�21O�AaRП�^w������H���	�Z�*�����"����P��O|q#1�O�t�'o��OR�Ưp�m�C�F0s�Q5(�D9|��ل?���'��(��'�������ug�aݹ�t��?<Y 7��l��ȁ�aӌ�	%�&�D�O�< S�?��I�|�S1��p��]�+�A��W�eЊ I`h��<Ѳ�ş��I��u��'��d�9^<��i*�$`JW)I5�Ira�Q (+�- $�@�6�p7�f�8b4��㦝�ٴP�Pպ�'������.$��t�c�ԷUJy0E�-h�l��s�������I��<��韐Γ\�<ϧ ̡`Uo�w�x$� C@�\P��[ڴ��q�����OP��Y�,G�+T�;6�b����%E,D��A��R!Hn��S�� qB�5��|���%��y��R���O@*��� UB�UC�`��_���`ι>�J>��T?ّK��"�p�瀭{HN��f�7�	S�}�'3v9A�ǉ28v�Rg���N�M�
�'�.��s5/�v5I�$��P!�'U�8���6`E�@�daC�e�p�'��!�I/~�y7"� Z+R\B�'�6�IL�(9\���fϭNrV��'�2!�B��:}_"V�C���[�<�7l��S�!2�ꃺ N6t���Y�<��˽\���P�O�0v:���_�<1@+V8P��i�M�<8 �Z�c�Z�<�lٹ|�lX����8zE8r�I�Q�'�B�'�b�'���?+� �E���١Q&�]Z6��ON�d�O����OP�d�O���O@����
����SF��btD5pѧB�)���oZ��@�	ş��	ɟ��IğT��ڟ��	\����Ȃ%Z[��q2j��|�4�rڴ�?����?���?���?���?�����2W�ʷ�����u^	zT�i���'���'�R�'w��'���'�
�F.ȓz�h��S�n\.�ѥ�fӲ���O6���O�d�O(�d�O����O�a�i�
L9��s�E�]���PCUʦ��	˟��	��	����֟4�	��RA.d�t��  �/8�Fx��J��MC��?)��?y���?����?A��?��,^�Z����2�,gU"%[1 (.����'��'o��'�B�'���'u�jՔ$�֔���6Ypj�Z�����7��O ��O�D�O>�d�O��d�O���Ԛk'`x��R	p����&��o����I�x�I��4�I՟p�I���2D)a
еy�H���DF�v�Qp޴�?����?���?����?����?Q��-#f���7|���+��F�eL���iY��'b��'.B�'���'���'#��xg&��j�,�BŊ,�Ŏ{�B��?!*O�#~Z�}ɾ�1`$?$\�8�ğ��Mã6��o�'F��;OJD��MU2
�`���&&l�z�'Yr2O.���r�P��ٴ�~"�@wІ�r6��%b����ׄ�?�'���䊽�hO�)s��B�-_6iu.}`�n������O�˓��lśv�C}ܓ�� v� u�(�@E јG4������g}r�'U1O:�'9�̽Cq�O�L�B�ҴN�,>0�'���V�O����O�)�-�?�a�����:RjT�si��5qX��ý<Y)OZ��x�UM�"DĠuJ! ������O6Yn������4�4-�3�E;�����ݟ1�еڳ$�O��D�O��d_1�7m??��O����n��{0M��G�4s��G�\4�1�� #ړ�?.O|b>�r�#O�F-B��D�6��a!3b�<	D�i�P�=����͛X��@D��B�a�lo��>����?�'�>�۲�7-��xB%A��cŖ���"�zlҒK*?A��F1L�������ē�T���)���IO (�$D۶23��������& ��<!d"�(0(&U"�=*��T+s#Y��<
ش��'����?����y�D�RCx��ߥk���H�hG�;/R�qٴ��٢=%N%1�Ot�O��M�'|�)i�!�v )��H&X7�O^�[���o^f�94��#`8�ň!�'�2�'`@7��̤|�#�ic1O"1AV?K��
�[:^Q��ן|��'���'�"�rG�i�i�Y
P�Tm���(A��MФq��ޅu�HI�I���'��	o�'l��l�7�@育��l���#��o|Ө��a��O����O��'<�����
H|�9g��2WU`��'���?A���S��*�f��qDG�.0�uE�6j��C�Lɿ�t�+�W���6$���LL�7�|���n�17�(܉ȭ[N45��I�M;��/
�@Q��c�?��M��k�+\�ъ(O�HoT�9���͟���N�b��h"���7tPE ��ӟl�����od~��ؼ%�Jx�����Z	��XF���Z�@����Q�P�l��՟���͟���ٟ�OEh���
��ڀ�L,eY�Lː�i�U��
+�'>���O�b�'�6-�O���p��'�`*c½WAL��*�r�'�')��''2�-5���6O�1T�V*V��+�c�?�>����Oje�c%<�~�|�]�������'������Sb�aJ���D� ˟��	�D��Y�Q��~y�d�Nّ������O�e���X�l�E%6���E�O˓�?�VV�<��]��G�j%�b�IU��l!�%Z�^`!��?q�.˶vj@@2�O����<�]:c��P���'4j`�ä�%���� �$8���'Jε�P���I<�,p� 74�	ӓ'V�"�@�X�0�n Ԩ<�e��2�|aF���<��F�P�BKv����NQ4������������0��E��#`p�BB��7e�r1:�KL���C�A!:���������̩0D<�+�S=w�2�I�	Դ2���y,uYe��!k`!	'Z+
&ZVDU�KBR�s��Vd����kQ|���3�AȆ!W1>u���CZn��<��ē9�0�cK�9}��@�͊)hpc�)	&��{c�Ix̀�
�F0�N�p��ɹ1k�� �MJ-�v�YweN�:li��@�+�H] �P�oc�1��,Ɲ<� �[2�
�&u��`b��(�M�������_�Sr�L[&�N�n����*ur���d̻v�d1�kӄݶ����GZ�К��+��m���2G�@�w"�K!J�@J��������1W�T
G�sy��'�B�'��'�R�'� M��]�b�]A�J��PP8y��Ӄ$u�'`�'G�^�����|�'�;�r�@�m!B^JŒ�*D��	Ο�Id�IΟ���v�(�aWF��n!���ğ
j5�'��'>�X���A{���'�X�b��N�oJ��@�MW�#���:�'���|�'�r�H�}�1O��Uhޢt�T���"
�`�t�J��'��'.��v�O*��'�T�ވC������?�� W�@�?��'B�'��MYf�'|ɧ�ā�
A����O�eoxL	��F�?,Odȕ�O����O��d�f�AI<lS�� k"���m-?��m����?	�M�fGx���@��(���kF�)��Œ3�ˠ�?)�;�?���?���:(O����O<P��
�p��̘��Q���O��i���O�O>���Fn@��#���u�<1w�Y#^����H�Iҟā�TGyr�'M�'=�D�#w�v��!�<���h�k g�O������O��D�O�����{���a��R�_����O��D��$�n��?y���?�L>q6.�D(��-���ȍ0�Ó��D	  6>�$�<A���?���\_ �dA��6Y�Rt�vJ|��ءB�<a��?	����?��=ąqN��Hr�����4��2CL@����?����?a(O�}j����?���Ga����� 6�lPu��Oz��?�H>���?Y�����y��"`�*�SoL%.@�b�ӫ���O�d�O��N��}�*����"	�ސ2�Dʧ��Bǜ8�����O�O����O�$���)� 4���� �l� �Z�2����O`��<�@o����i�O���ퟀ�(VI�հ�;��u�p5��=�$�Or��I�k������Y젹�!�*n_&���� ����<�� ��?����?����"-O�8*�. Gm��6�T�tQ �f�O�$�O�u��a0�)_�H���H
�4�����2�?���E����'�"�'f��N=�4�N@B��ְB=N��5��3�^t+�I�O�����Of���O����L��<A��JbP��,�59�t���KV���i�2�'r��O�Yj�O�)�O���=� �3�mO(��3I�t�J��'���'���U��ON��O�)2fA�,gf���BR��`�����OR��H�o%��&������Ily�jG����ܫ[����7"Q���Ip�Ο��	pyr
h��:�F�<u�(��+�e�q��!���OH�d�O ˓�?)�N�l�i�.Jqv�y�E��(1��{p���?�M>���?�-Oν2���?5�eކl���*"e�p=��0�<���?)���d�O��D�6=���[BZ�k1��&�����Ɋ;l����?a��?Y+Op�C��j�S
�1H���g/���ck�6Q��(�Iӟ���\y��'L"�e]b_>9�T��_�Z (`.Ԅ�Y ��ɟ���˟H�'�#�7��O��ݬc��FF�,H����"V�:_��D�<��?��M���?	H~"�wr��HC�d�J��FT�<^t������=\umZj���'��dī<��oَE�Hb�!w���`�,�������Ls� T,&?��I��R͠��D��?n>��f��
::�OћL��',��'���Q��'f���-U�jJ�g�!x��8�M_�YP�O�r�S�O���h�KL7%���fL��#tl���'���'����)
�O6 ��*�1��	R"ӭd+J��-��' �ͩ���O�扯M�Сk�h&�<U�VC�-[w��$�O��A��<9/�|㟤C�E��#�$�5 }��D�|y��ʚ�*���y"�'����D�"�BjJ��	wK�%ylҹ�%�� &<��'�"�'��OF���O��c�L^�TC���`��!*�$L郬9������Onʓ�?1� �0��4h˸A섃�l��HD�`΍�?����?1���'gB(�@����ɔ#�8ur6�P�Z��	*�.� yN�'�]�D�ɑn5~�OTb�Q:S<�}Iӊ� �\L�L��b�����O��*�X��OfX�h�*4*��ے~�Pp�B�'��P���	�4P0�O���'���C/�^C�NPb%3�C�h��'c�_�ā��&�Gy�]���	�xĪRKy�Ka�ԗ'�V8�Geӌ�'�?���K)�	��N��J�`S��ED��,���O����9_�d'���F˧e8e���;9�:�R��O �!q�W�v�K�i��'
��O!�O�iCR�x����1u�H�D�����$�vN���Ov���O|�)�|�'r�}�s%C�<ɐ�R�[�>���3�z���O��d�<;q�U'��꟤�Ɂ@GL�Z��W) �ī~a��៼�I�<�u)�k��Ob���OZq0�E{�1���0_�u����O��$�4c�'��֟��ay�m$K�~P:g#�(e�r��PE�>@`b�'8���'�'~�I��,�����'S(��v���|�,8�k��aeZc@�ko�O���O��d�<���?���D�4r$��\�S���ȡ�ַz�Q8���$�O��$�O����Oȱ�QmXަ�S>��Q����F:8�h"�ş�Iǟ���ȟX�I_yB�'��ڜ�M*�OTȜ�%ӁD
F��O���O��$�O�\Ѹm�CP?=̻W�D�a�(��(s�O�aZ���ǟ��'���'����y"���ڢ"Ԥ����-	@z�Q���O����O�����HY?��	ϟ0�S,Z�`T��k�Xĉ�$��P�'��'5�A��y��'r���|� )��h3��/4 �g�ftd��KyҦo�V6M�ON�D�O��IJ}�[�d�(�H�5Y�@��d��4�r�'�ҨW��O^c>���+��6�rAs��q� ,
�O�qY'M�����	Ɵ��	�?���O ʓ�Ό��h�)%�xz�Cсr��x��vgDΓ�?9/O �?��I���H".F�X v���M�u�h�ش�?����?q����r���?Q���?���7�*�¢e>TR\��v���{x^�	���?I-Oȵ��!<�	�O����O�xz"Ř�!(mK�l��m$�upG��O��E�7�vtl�����$�Ɋ���{���NN�
��m+g��(���<�g��<����?A���?���?��K���w+��p��"M�: (��� ΁����'���'v���~J*O��dM$��xr�^f��d!��R�|�?O����O\���O�d�|Z���+D�v%��^`�1!�9ȴ������'��'���'��I֟$�$�d>y�4�e@�C�x�H��u^dy�'U��'���'����PH~�Z��O��a���y�tT�2j�6nv�C��O�D�O����<A��3���'�?!�'ǦaR��
Pyj��!�������?������B�*�D��O7r�'���%0$����&���В
�� ���ԟ@�	�t{V� �(On��*�5CɁ�qt^��Tc�5t�>�$�<Q�;՛�'���'���Ⱥ>I���#t=�� ��<�Zy�
�>�?I���?!���<1-��d/��J��TkB(0�X�#fC=zO������n۟L�	�������d�<��F p�t�����%N�闬���?QBB��<�I>��D�'�^���M�<�u6#G�e2�8(��u�����Od��QD���'<������9`D�%�BV�&�<����j�Q�	ҟ0�'��XE����'�2�PI��LГV���c@�K,��`��'�b��������O�˓�y�bũ �l�@��|�|��U(���Ę��O���O����Oh˓NY֙q��^�*�[�Ȥ���ISy��'%�	ӟ���Ɵ�� \lQT`�zD�Z*v(Z�Ea���y��'#�'8�'�	��v���OȺP�4��BzB% ���DY�	wy��'!�I����Iڟ�@�`�?mk��Hh�� �ˢ5�H�[���O<���O��D�O<�t:!��X?Y�ɇ�%z�$�s��xq"�K B:��	��ܖ' �'����yrP>�� ��zl�)�!��!e���@��8�	�H�'RPk�̾~���?a�'��L �MT
+������A4�Zɩ-O���O��d=a(1���v>y*�+.I0��̑g茰Z���O �$�O�`A"��릅�	ƟD���?U�蟸��y�����E
���:����'�ϗ
{�|�O�SI�=���Y<o�d�G���T��G>I��xlٟ��I��ӧ����<)'�^5>����a��'
�PG+ƞ�?��$�<9*O���/����mD�3Je�
��M"Lx��P�MS���?Y��W��9
7W�d�'�"?O�0�`�����ĩS�tM�����'�"�'�b�d��O���'�rKST:��r5��	�PM�C厴��'��e�pbuӪ�$�Ov���On��O��8(�(�
ӗn
��Pdɖ1o��.[�&�?��?Q��?a�~� l�"��/<DD���J1B4�!�v�RW�V�'���'��+�~�+Ot����2�1�[������u	�3O��d�O��d�OV�Ĭ|d�� s@����J� �:	�p�i�i(������֟�������'[rj����D� L��T`��ڕ-��E�d*�b��'Pr�'�R�'�R\�(A�7��O��$�T�liƇ\.�X<�!'G�J@����O����O���?y�]�|:��y�m���!L��TP�#�?y���?���?qQ���ƛV�'+�'�����:O�61�4��9�`����u�b�'l��۟��&��e��|�ņ���(*�+�T1е"2���?Q��?ir�ͩ_p��'��'��t�O�ZYd6m��eԄd�$:�bX�-���'!�ULb�|�OL��.���l	]�N��bFH6
�n�D��y��l���I̟���"���?y֋�%^�h�A�o���KA@�?I�@��?�N>E���')�SD`��n�Š����s�|�:3�q�"�d�O��$m�0�>���ybbE�WB��y�aF`���1E��?YM>�� �<q-O����O��T`���b�J:�Xt)c��6sR���O��%��W�Iߟ��	q�	P��(q�Q���@�[�D��ݔ'��aP�'N�Iʟ���<�'�|܂��ߥP]�ղ��������O@�$�O(�OB��Oz4�n�a���#wŏ(R~�dq�B�x���<9��?�������&5����S�s6![�Ѧj��k�	��ʓ�?�����?���Z�*8��L]6`���Y�Y�T�቏�!���k)Ol���O����<y��/e��O�Ir��il���K�>�À�'�B�|��'�r��a?����..��ݻ�&�Q�tz��ON�$�O`ʓl2�郛�T�'E�T�Xjj|��a#Än����6`�k�'�"�'��1�'7ɧ�dJ�Sp&���FY#*�YH��A��?9-OZ��Ʀ�O�O�6ʓ��9H5�v 01�d�cYV��ß4�I��#<���S�\ ��`i�x�HS#��?��.U��&�'h��'|�$�2�I"���Qf���%'ȹ"����g�O�0��IA���?A�)�y	����N�
�&��c@����'��'��9�-3�d�O��y���@l��(�6-�S�����G�O��O�ɠQ 9�i�O����O���F��_���th�Jƌ{c@�O\��P$��0%���I��%���'Z/�B�ig-�rҮ5q���pyrD���y�T����ן�$?� 5�ɠ]���eO�<��2p�۲;w���M<9��?YK>1���?�M�W�v����O	"Þ<#f�%K�|��my"�'�����$�O~������CW!KFҠ�cK�>G��ğ���i��ğ��	v�����	4m3k� df��:bd�P� x�'��'��]��A4΋�ħo��CuX7yځ0­OL�(a���?�K>i��?9�P�<��O.<9��'RҐ�7䄣����@�'\"�'B�ɗ+�Z$*L|�����sIT�g u�5oU�lk��t�^����?����`��Oh�p����~�B�:N�!J~�����򤉃C>%m�H���'��tG�<!�I�)����$���D�����G�Yy�S�P��\�S��� ��u��=XYʰ3b��f�B�Ux.6��OD���Oz�	E�i>�Q 
<�d,*��ȴߵXN�ʓ�?�/O��}:��u�z��@ݖg�e�E��rJ:Ͳ�iU��'����\^�O�)#?�-WG�@@�.ʰGLpb��^ӟؗ'�� F>eV�O���'GRK��w��@b��Ѳ<H*��W���mf��'��9��U���O���|���|�^,H0�̣�2� ��M�W�	wp�0#l'?���?����?��@����Y�Oe�z�e߅/}��&j�}	���'��'S�-�~�<qƄE�-~�@�~�{��&LCH>1��?����?)��E�r�q���>=(@� p�]	Ï	U������?��?�M>���?Y�ȓ�/^����ޖ$u��7��#sڤ)���7��$�O����O��OH��F��|"�% <�Q�3(H���lX����?aI>���?�%eC7 �E�O� �H��Ã�l�����b 3lR�#d�'&��'*��'@U��cӂ��O�D�2�2faR�+$��B�cA/h<:)�S��O$�����e�O�p�u�R<�E͎��4���'���'�:��'�2�'��O�B;kg��-fhT12%Z�2���
��''r�'�̤�q%ߘ��O��l�� x6\�c`�1���z��) ��?	(O����O����<�oc3&�Rǜ�V:t�gl�"7anʉ#�2t��y���O:$��D�l[*̲d�U�x�3���9��ǟ��	�����ßP�	�@�	؟8�C�NKy���M�=�����V�u���J>���?9����;w�=uExiP�ą#Q�u�)O����O����<y���s�X��D̫X��8�g*ܾ!K.��/O��@�I�0��ȟ�	���k�e|�6uX��#?�,�`�ER> ���'���'���|��'��NQ"!^$@��=/X2��0��
-����ݛ����O��D�O��$�O>8i�ߦ�r1 H<>h�iֆD5eȁ��Ƛ�	�T��ԟ��?��%�y�H��� �[��|�层'���D�O����O���O^�(G(�|J�!�(�ś����"��"e��*���?I>!��?)���n���OV����#$t��a��'���f�'�2U���I�B�u�O��'5��HluԨXզԁS���q"@��'�2P�(�T�*:+<m#U&�� ���UK�!j����DJF^ m�J�$�'���o�<�qC?,�@��+օ�=Ӡ(���	ܟ���=�S�'K# ,B$m[!r���G�-:�����
>V�M9�4�?���?1��U$�'�r��>7/j`*4��^����G�.D����'=�-�z��HH��üR�"��D�q���d�O���<�x=&�$��㟰ΓK����R�M�fG�lA�%�%Pg\��?�#��d��?	���?�aA��l粤A��R{""�Pۓ�?��
i"qR���'u�Q��̻[���V��#\̍jqk B���	ʟ�J3�t�$�'���'��P�aW��qR��s&G�{�
�P5�H$L3?��ķ<�������OB�$�O$!VO+�6=���Z�QQj�C�f]G��$�<y���?����$�$Gg(��Epp3A�$��	�vD/���d�<�����D�Oh�D�O@ s>O`T�QF��gtE����s ����<��?������K�{$���ON2��<=�a� /V���X%��'�I�p�Iן��s�$�'Ī�+wς��MⰭ?��0��?a����d��i���O��'��T�L��IZ@烡J���?{��Iݟ��Ɵ8��	|���IAy"=��B�ڵ��t��!:@Ќ���'��I=J��[۴�?���?���h�I5R�z	goEn��3���9Ψ��ПP�I%9��	j�I|�'S$<|{��Jm#r��#1
�Ɯ��6[������I���SDyR\>}�pLH4x��1�p��}`$qۀ"�����Ʈмs�"b�"|��dF��ȣaċBr^|���{}P�P�i:B�'}��Q+d�O�i�O��dG�8�v����5-�� �#�"%���T�5"3�˟<�����/ 7I� z"/,H�l��`&��|�	+w���'��S��&�t#wfƙ]F��+�.O���ܫ �Gjy"7��8�ON���O��ľ<���]QZ]���P{L�pW�۟p3�"�x��'�2�|��'�"��%���Y��&"�4�Ȑ�j}<�J�y��'c��'Y�I?o��U���"=�����X�U	+HF�%����o�Iߟ���w��I�c_��S"]!��홲��%1��O�cE�=Haje�����v�\�$��57EX�s��UVـ���ǰ�Ԅp�����lq���ϟ|��X�IԟF �	x`*��O�D*䟈��I� O�Y�b,@�=���`��O����O�O��d8���1P�.1D�0lڑ^�����OP�c�|�6�U7i%��ȓ!T��+\Z�N�f)Ш�xp��I'<�ꍀg,R"U���Ă�xD�Q)#O��'f�̲f���V�i� �,����#�'}�2��U���l��i�M��>X�s䮝�b��ɺ��0XJ6)B#�Y��+B��ԀB ӯz�ZPp��k�x�� H�'�
��D�8e$-%I�6��D�!&�5Nyzxt 2�MKt �!2�6ٚ���Oj�y ��OX�d�OzMq��O
c�֝����-�6\
A��)X*%�f#?�rFp�OѤ�Sf��8��_5]����D2x��'��O�M�6i��C�8CB�D�<q[�O�0�)�'B��L�$/ũxt�)�ޛd���ɾ�~rȪ�TtC f�8�1`Ϧ"��ʓ)�*	�T�i}��'	�P��IӦ�X�aD�6�����'$��1���?�nT�3�2�(͎q`�)����))�i��!A��0˸=�Ç�h5��=8uz�9�\=v��ʢO�Z�O�<p7I�e��zb+�X�,�O� ���'�┟�i?�S���1�f\�^ѶQ����b���'���'�2d�$��1LoA�rGΛ9IxI���Ĝi�O������'V^�I�둭����d��<��ʈj�'�?����?Y��<���z�B��&�F�)�QK��ACJ�5�(}�`���ػ�-&���Z1 }��UG��[�*�`�P?b�'�p�¢�4���O� Diق�E.7aj�Q�P7�0Q�x�#�=�?	�COj�$�q�x�yv@ׇaߒ	�ȓ{]Ry
�ܔ+�����]H{�����"|�"e�FQ�����޼E9z�� LM0�4�s�/�?����?Q�FP��Oz��`>�!
}�.\s�bW<|������iW�q��'�F��4�t�yw�N�G���0�V�g���	=b�7튠`���g0�������/��<���NܺU/D�=�<B�IV�s��x���􀙧O_*nj�qj-�V��O�)�>1�V*r˛��'�B�i2"�)q�S��\|x�U��%#�O�h @��O����O"�P�́7��ybIUc��)�i�=�sB^�W�WbK�i���Y��&�0�,[�`ԣ!{J�z��B�����������T�ur C$O8P"?IS�����~�R��*�Ȍ���A;ǰ�U!�D�<i�i�(aRi��g�>_�P�Bf��P�'hB%	>��X&��>�̨L�pj��M����?)��h0��Or6�����:!�۶)�v=z�f�,S����	�1t��mW�tOvX/���|rL|R��:���MY�=���IPnVM}��^���9�I@Ҳ��0��q�8i�Q��WP�<p4n�,� �z$q��쟔�����D��bϣ1�J�����5Fs"��O�)��Iǟ��I ����E��d��4����br.�>���S[���	��B78�tt� ���$���?���eQ 1;6H��?���?������v�Vd�B��,�Y���G� �P�"����IASrA������g�/HT@�+���Y�7fI�p����D	]}"*ϧK���3��$�o_�� �d��?I�&�,��'x� �ɰ<a���t�B�+^��J3z�<�A%�7�v��u �3Z�HQw?�C�)§B�r�`���_�����	({\i�!�-�������?����?q���t��O�� H
RFhʐ*6�4�#�սN���H��B��~�"^%/`��5wc�p�q�F�L��e�5N�@���C# bӾ���� ,���G��%0�X������t$������4�?�����ə����f��a�&���B�	6+!\���I���}cV*?Mx�'�ꓺ�D��W-�!l����ݦe�%�Ґb��ث���/��E�KT&�?Iǈ	��?���?�e��E�|���|ZwȞ	���:#5X:�I�9`ة��$ �:6�Ѩ1�>�>OLL\Hb!�� oV���K�A
H#?ir��T�	��	�;�&�D&<{@�;w�Niրh?�����h���38l:,�C��S�H�eP �'���	�PaH9x��GF�䤰t��q��0)O�����Ŧ�����ĔO�>����'���,Z 
y��!1���'�� ,�b���(w� X�ʑ�i���������'��'8."x��D/4�q���	4���'4�ȸ�F�HN�EitJ��ȟ��X�+�JDZ����q�JL)�$[y}B�2�?A��?Y��H�Ju�EZ��Nѕ<KLqS��>!����=1큶4[<D1VA�p���b]j�'.�#=y^w���� Ɇ�_��!ڦ��hRā�'E�'(ay�M�^�2��f��gk�9��.T�yR)\�^�(X��H
`�0���nգE��Y�uhCN��Lx��'�J�m��'��a�'��N�@��'@�ę�MҞ�����'5��y��'X:p�bL�F?H�R�*�0 6�0��ia�yIF�����aKS,��-��_f��4�F �b�`O�7���ȓ���(ǎ�`�|a���S U��8��(HR]��JB�r�=
	��\�܄ȓf3J��(KU��I5HPj)n��ȓ	#
���[�1�4%�(�:#�Q�ȓ"�æ!J�2����ĄчȓpE�b�A�<3�-�$��%b�ȓ
4�� ��|�x�BE��z#ֱ��9�v��H�����WjR�#\�Q���Z���ޡ�qS �]|�q��?⾕ˀ�N�M���j�t�@�ȓ���
@Dz7$���n1��(6��zB��&X��,����6Lh��ȓc��&��l�ѣq�L,7�ԅ�S�? B���'�B.���G5�b(��"O��� ��Z��h�MMy�$X1"Oh4:C�K4d��8�MYf|R@kV��(KQ�#���$�"|r6/�/=
�k���~
�H9��~�<1��\&U�a�R�H���{�i�9/�(�����f����gܓG����$G�����Ǣzn����`�2�ӥfOI��a��H�*�2"GʶYmh�ĄJ^�����*�[�ꍻ�J؁t]���.�Tup���/]�P���J?)�!ʉ9]mZ�Y�*��H��y�t�:D� "��ͨt������t�ti�@-�>A��� �k�k�a��e�>o��y!�
�0�"%�6̛�ybiܚT��!s0N�1�*W�Y�̥mZ�d�aa&֠E�2ţ�����,扉D?V�Ț18��A�pÚ�g����L��f��qiI^���1�ʍYUFi�#CA���\�L�"��T�e�93ay��K�tt`�e�U�R�t�Ñ��O&�#C�,~�.��7t�|K���`��TBc�WwOn��a&�-�����	e<)��i���B����jC��� Z���D�? �I#����lY
�E�l5�S �5��
�$�6JN�h#и�G�/"��ȓ9��� �ER;� {s�O�[؉��Px���147����@�\�S�63�-O�(Q�,ω!p����A�g):GO� A�lϦaG,�g��hP���/�`
V��4�06H� �A�"Of�'�ڌƀóv���!�E�i]�|H�C_�$��ŏ��ΨC��Q�b,i�A��W��f��q��%0�i&�OnТ'�W'�z%�"�����Pe��B$~#XE���_�Zb����ˡsI.�O��̱�G,,B��� <G>�A�}��N~Ԑ2"�S�Z��	� K�Z��6�&?kpEH���X�(=�d��iU�x�f7�'�~r���] ��W&�˅ub������*�O�x��Y�쳰C�j��ks�ƖP�X��'ֿ
;M�f@_?3�tTa���||hםN�'�H�Y�?�&�*�(л�@�{7���#��caQ��"VF�>��%�Ȇ~�,J�Bѭ)�8Lʕ���xy��y�#6)�F}BC�X���7g��%re4R0D`{�(�%b��A���'��u��'FH�R�xA�ءX���[ �~�A�74�d�S;��8��H̓R>��XvF�g
lc��	D�|��*WI��!��:�b܊^H�Z@�\.w�l9BbЫ)Ρ�e�o?���N�����7,ݶ.����GNN����������䓟:>�u�t�r��M���"j=�>=qG�-���1AĞ-�����(���{2g�&D#���5K0��P�M<\d� V޴�mq�D�:����5&�A�'[
 c�Z�w΢�)���0��o[[8�Qa�%v���aa�C�X����`d���:�����Q>��%�O��U��O�!d��=�Q&����1R�"�6DO���pE��GϘ�[��P�sI�$�- X�H@�&D^�|6If_��q˙�jێ�3&B�2��TA���ʰ��K�	��A-(h�ZP�̻D*ɋ�Q	n�����O?��<V"l��5CFC�E�%��L,�Kub�?]3n\q�A�&^���D�~�aቊv�|C��ӫ�ӂ��%����tZ�!��a_z�!�D�z5���g}�@*�7��N�h�p�;tڬ���^T���ɤ��ԴS��I��ܬ�-O'C[pb˼>s:�S���0qMP�9CKP0&���c�:gz��I�X��Hq�_�<�!�}P,�j�py�0eUF�vH��k�u�'����]�.H�~r���*$R(ԁ(8��B�O����2�RBD�RE�Sj��?!BR� +?��'~�D��ѻ+ĲL[ F�?+41k�'��Y)�E�B�S�����%�B�V��H�e	�($��҆nK��y�L� e8x��+o��x��ޜf��x)�e�  ��[b��6�hO����'�!7T�`��'�A��?yt���'D�ZD3$�Ü]E@� �8xC��D��R>��Z��\:�"�Q�E�Tb��z  Ke?����+��Rc5MT�`3s�>u�����P:���Dr�	a�Q7G>-�U�P�E4V��45I#�R�Z�rdS���� ���&��A`��)�,�孊=[tkbe2�Od[�%�:��Î��׀�iQ�/y���"����x���8=����"�Sm��PvM˲�hO �Ȏg��@��$X�;��4����=K3�+UB�8�y"e8'������7A(jU�R��ybB�
8%"�j�O���K¦��#���?zu�ңtS�4bе
*°�v��l�p����2�y�_D����#�b �ŏX���-a$)˰[8(Ј���O���WF���	B
f(��Ͽ���e�F��炑�r)b �ū Q�<b��R�])L��l��U��!�v�(qߕC��P� /?]���'P�Et�.�ɯ))��"�!]�|L~����=pN����-W���c�"זdf�B�>[y���'�<��Ap@+W�*p:��=yzR��S�? �I�V�_�� ��������?L���틾+>Q[t�V�N4�����T�Ӫ0�oET���+���wݘM�r0D�0J�O�1o�AA"���X�H% A��#v� `a3��!�T��e*Ԃ�>27�3mq��͒a�L���ޢT��pА#ـB�!�$Ύ&cНÁ �;q�~<ʗ��7z���P�Ɯ��c�G�z�"P��8�ԉ�!��8��'��ɡA�*�����5b��2�D�1;f��#~��X�@ d_�P*ƌZ�h��"���0FP�%�gƼ�a��&\O��Ƥ)5
�[#fN� |���b�	�YZ Z�M	Qm����7�8���!wܘ�a$�S3<u�H@�ɭ-�м��:D�����"s�� r�n�+K�����/ղ8� e�|���$	�l����RK��Of���\U�=Їe�Ύ�i�$�4A�!��Y99p:k��\�$��=Y%�"����G0T���a��[�TSy R�����$L���'���谯^;�h*4��<H�j���L�j�ʧ�Y�2����XX$����}�r�b���Uj�:
�4����'| ���8*jJ4�#�-.�%��}��K
nŲh�qd>#ᬠ9��<�������?y)�k )\��h
��.:dx0,&D� �G��t-�3B�
o�T�H ��!{�����W�>!���6�� �B(�'a�L�'h+�nۊLO�D	�i�I�QEY*m.!��*)7����K�.��1���F����>	�	�⪘3YF�t�P��� �,��',�I�VN�-mڄ����<&���xۓ����g$��R����l���`��Wn�MKH����f�;=©%&5Fr�{���.0���d��>b0�3�B;��'g�X����g��@�#��5`��ͷ�Ji�:�4as��#L��0�q�!@΄B� ��� b�GY9�S���L�& а�	&n���#_�b�e�T����~��w:X��FW���gj��qQ����'�^=@G,F ������� ��`K�+�B|�Zd 	�}E|�X����� ǬD�O}��D:2	�E�Eo�,�J1�b�i���XgfA�	�џ��'�@���ţw���i��3��Д~��`��߸
����h��!�E��d�|��t1�l_8�y�$%�������a��LY��3�HO�%p2��K��p��/^�C|�$�Q��?Y8�dO:����� m�B0�C:� l�N,�q�Z�PN��E�4kś9h�)-�3XL|�*Ο�9�G�'ڒ$�e�����D�ܴ^���30�À��4�`/nԬ�E�?�6h(O(�a3�3?���G��]�Љ��7���"����~­҇MK��ed�!MF|`D"	B�~��lç�l|15)jA���{��\�g�̝n����T���J��äK�(X�31Ҭyj�_������n�"��'���H��G�t
�kUU�@�F�B�+������.�'o�D\hԇ�Z���!�F[���P�<1��ۉ��`������h���;� H�0�Q�$m"Ё�`��6"=<O�ъ70H�\�C��I�� 36	��]+4P3ä�<���f�����eM��� �J�RFD�" -VT�!�ʗ����D�c�(pE��&��t��_D�F�+|O��P�&�$xMt �C�,��E*D�'D������f�U�6t�s�b͜3�fT:���7a\x��I���u¶��1�ʮZ�ȝ�>���-s% z���W^�P�wj�{s0!b*ſ,!�$�%	Ѭq�c�7����V�!���<򌂖��/9(�����!�*v�>���$�;ѹ��6L]!�D֗̸�©�0ڰX�FϦF!�$15���� L^�d��|x�䖒
�bG{���'�2�17o>Z������)��3�'�r�B�����8����q��% �'Va�N
$
�J����V�D�Y�J��p>M<y�g�{�@QDMP�rڊ�`���s�<��K�z�89�Ђ̏d����o�'0ў�'pL@)�a �-ov��c� ~54��ȓG��T+B�gT���D��]`@�x��)���`�$`�2��� A�f�hwG"D�蘧�.kX�]�/��a��)6���\����<]V�h4��I:�`�mU�r�H���=���b��h
�n
53��0!�Z�C!�$�]�0M�f_`"(1��HI�4!��\9zHE�%�!b�)�6'J>!�D:MFXXri͌vD(���S$ �!�� �h��D�JE�Zro�<S�Y	A"O\��CI&6��8�S#Ӟ=r-�"O������x%y���
bv��Ht"O�5YG���)�`�hkVт�"O�8)�FB�y����q��&?U���"O��F���HH�"M�%U@9��"O�ف��C1��uZ��ύ�ZLi�"O.u2�ר3��),�+(!��:完i�k�9 ��BL>q�!�d�b"��,��j��r�!��ݙF� ��Fl<.�h���<t�!򄚲r@pĊE�S�-���P�ǝ6fh!��#@ld���/�4ie�(b!����!�$��d�R a�?	Y(�#�}�!�d1z���)Թv4��!R�!���65�$Zg���t���]��!�Ѡu0�SgE1�)��Q&!��R�M�.����W e��@��$7d!�^�<�Ҥ[ԯ��j<B���X}e!򤒚�^�!�"K!/#�2D/H=O^!��XC<ѫ�[O���uI�dE!��F�b4���f�;:�}�dn��b9!�D�Q��}�ҬL?-t�
,X�T'!�=(E"8�`�],2��!�Ě.qB��G
4f����՚.�!��cl\�a���"��ɥ���<j!�ă/ 4��!:�(@	�
ߍ%<!�$����lǽ�0Hc�+({!��:7
j��tP0�ܐ�FL��3Z!�.ax��d�̍e�fm�f�[CJ!�RCarq;�G���.pAC�!�!򄇤:��$H�Mut	2Ta�4>!�����4�"d�9R�4mʣ[�]!!��H.p���s�مHԬ��e %f;!��>}�]����!\�(�� ��)!�$��]�ڜ� l��nŘ��&N�!��k��[��  ���!�q�!��.V P"��e �$��H$7�!�$To��A�D^��̹sk��B"O��
�L�_^� ���j�j؆"OL�R��>��e��e��1�6Xx�"O��S��l��04	_7z^���"O��2�*,Kͼ��G.T�zW�x��"OT��'�:#�`�/�"1�� �"O�}A��қyδ�R�)܈#"O��gE�O�< ��Ԫ(�S�"O�5$�� RМ!��A9���Ѣ"O`0�B8[�<� ������"O�cu���"ݺ���n(X�"O4yP�U��K��G�
�(�!ãR�R})uL@9#q`���*\j�Qf���
h�0K�'�4!�dԲ>���@O�cSN��cgB�32!�̖L,�I#1�r"����H&z!�X_�l�����T:P�P��B�!�����M��fH�	��?�!�$��N�6�5L�e�p�CD��z�!�/w�}�UK�+���0E	�~�!���?qV��rčQ)	�|��䑮Y�!�J�S�v��r��M~�� ^|�ݐ�'�Nh��H,NQ�A����ob�IR
�'��p�Ŋ��0�B��"�p�0
�'oީ�M߲L�L`�Ҷ	BZ�9�'��ݑ�`��J���R��\�O��R
�'���< Ш;@g�
E~d
��� 8E �n�2%P���ߪwm�%r"O$�á&�?A�2��H]F칊�"O�ȐQc��#
���@G��aEl�f"O��1��{�0��"F�i�����"O��yAO��Os!d$� }�z�y�"O0*4$��U�jT�A��b�h�"Oj�(t�SJd�U�f!K��|)�"Oܰ�n
�$p��ru��鰸�E"O�A÷\_R�Q B,>��G"O�E�sk�1n�(�棒�8.�%�"O��۶!/<l��$��&r��ՙ�"O�)�p!�AB�j�nLpx���'"O�H��E��.R0�!��2hyb�!t"OjdI#Q!c����DU;k�@є�xb���l��ك��'I`%(`�S�����+��u8С��`L�n�VC�	�Q�Ni�AD���l��1�_�(9xZ��[�D��cǖ�^;�D���|2E^�$��d(J�\�xq��6�Px��n���l t��Ѓ���/U�m�&oA�I�P Ó@�}��g9��곁��g�$��6��=h7�%�C'6O��Ѱoʦv���(�;�m"Fv�ꘪ���.f�BI�B	��HOH}
� �:�LTi�h)���Z�\� ���R���3�h��A9N���#5}bl�.!b�8C�VD��@�EBA;��R2 ׉7�z��,h�׋�d}ʁ(�T���o-��x�J����3�b>�#?q��R�!�L�+2�EcHex�-�;Ct8�&�Ԝb�xaR0�U�c��sćBo�'@�J�K��!Q29XQ�V)-��P1��D<���W |��5�-��c`k9
)83A'��X[����2�Rrb�^��bɂ$�C'R�Լ��J�6:P�a�vԽ��B�v�P�cS"�����������1"�\�d�R��D�:/�a��W!�z��^62�	�[8�q��S*E9�����ΓO�� ��S��кa��=7:�P�[���� ລ��Ov��@�$(J�ym ��	;�)��Ҧ��V噇M��]&��9�Ӂb����[�/�}�%��3�0*2�1!˼D�6R�$D}C@��E���*S��HɃ@T�)�%�bA�?i�0Q���|�D���>v,$����)ډnH�8;���>9�i�"�脀 ���	�j�R��&�6�P�2�7z��`�
�4Z@	A���O���ӑP�F%�4�T�oR���0�؞t<y���+���aF����7'#}h�CT�-�ġ���$���Ɣj�Aa$����'��D�� � ���*Z��m��tQ�&(��e�����^�%Q���D� �*��Z���{����Tj�Od-�Mz�������z_"�1�A���AC�-��-��袏>��M@�Z]�ܴȐ�'�YK���Bc@=V�(( uj�d��cȱm��!eퟠFH��#�	�\ٖܙ�L(\� |���_�v��e�'�B�`�咴+���D�;n�vH��a��&�V�Ke.�&d|t���a�/��)�������'td���ă
�t��+L�ux�҄��#�a{2΀+_�����J�G��pçS�Bh
��S//:|щ'�$��^u�6��>�� ����	/.x�`0�#�Ug�bP�)������Ql�4�6�(���$�V�[�Q):��] �f��1L�
�-[zb��ϕ.%�ܡh��Y!r��ܰ��Ot(K�|�8=.�O�=�B�Q>�)���-�dA�K�*��Y�닒8��ڶ@$Z2�<�F��ا�H5^��! @$ ��@:�[e~B"���{b덅F����d�ف@���M�6�x*�X�
ވ=�>9��"�X�S��Phų.�����O9���+��K����X��p򳈐�\]4�X]�lY�a�';�y��ԇ ��t���3:2�I5��6�j�s�B���-���X�*��Q�����'�(=�B?�raKK&?�n1�咽.����*�PH�D���3C����9�� �-��17��'l���Q�����xBG�/�8H ŎJ��􉮰�I!?�J�a��	hҀ����d�e�˯4���#�)7W0�6�Zd?Q�';q���Ur�'0̤���LR�����+H�9ȑ+�<I��2/ ��(WΟ ��ҝP�.�'C�bC�i{��#��)a�ɹ6({x8��1Ϟ|��@ޕ��'��PZ�]�OTN��B�U�.^
-
ş���啮(�L��������Б�������a�D"T�$���&��%3��#�$	<P�$1���
�B�D{B�Y�A>L������$� Q$�t��Oh��P��-��=�|�C���2�z~fR����*�8�"ÏQ"K�4���oVE����6�	'��0��1}��j �M,`�V��',�(t dBƾ+����'�` C�S��\G��0>��n�@3�߾g��x[��䉚u^�,m� tr�+�9|���'��6m�*�@����6���E'ܪ,��!�6�ɿ���y�o�0+��X��i�y`cB�P��^?o�D��F =�ؙ���jn���s�^�?�`��+�?�fF��?����|�	��&N��!D��/��$H �x�K���K�H�/r^à��	:���<$N��V�duЧ�O#I�\�e�b��<�?�e��
8���D/2:�Qv���&ޭ�'&� \%� ��KNЩѷd�;c��E�M"Ș���:=�V�� F*q���t�Q&MRQo�w�� �����`<4��]}��r��',�	r�R9u�(��?��!�{���z)��J;g$,���ͬz�8�J%���^젵qbH�"|I�ͨc�S˦�V��2F�T>�Pߴh#|��T�Ry�1���?G�2ʗl�@�)�O	s�S�ԏ�{��50��w�DL�&"{��E���/.�����DԔ�?��*]6Yu�:��$*%;$�D���n�O��~��9�\�<�|ݫM�,�w(	�,����Sc`�`bק-��	S<T9�卨 �ӲF�H��'N�p{'"�"ݖ4��HP*W�L�R�!�v���h��۷,!����Y���Pk�'ޯF�|��'r�I�������4�q��Fd��O� k �T9n���E^I4p���O/ޘr���N6�p��ł����'�����k_�yp��)D@�DJ�LY�A�?��O˻��)��`	����0�8P�G1	)�a��
�:���;wO8Q	�o�?L��CFT����'��� ��`�MK�G^���A�;����?9vaϪlA��	�S�8Mt���U�d	��^��k�c̿(Ȯ��o��N۞����Y2x��&�-g�6��<_��!�WM���8w�-j0��1�;WkP@*��4?)g
%6.֡�P��Xg��A�t��?�cm��rڼ��瀘"��j�-'D��YWbm)�bF�
'f(jȋ
c�ԭ)��_8o�4�rF�T>�R�,�7UF>��l�j��/H�>���x�%Rv�C�	�,0j�#f��O���M%k����B�-}�ɋ 
V��	����4D,���ᐡ��'0 �P��4m�8���H3>4ÓZL�h�©��>�*���L� LZ��B`���TT�n�P���\�%o>" �)�@��
ߓ{�$�coȎ�>��V�J����'�4|��Z���u���y��ۍ{���rAz����B�s��=5��ȓ/��<�!��/^�r����S$�4�vcڣ]��<3��H�S��H�o'H�k�w�|8q��1m��Is�	{�l��	�'��}:�M�؊ݳƤJ".�J|Y�����I��p���
1/���t
K�;V��H �+�nu�����9"�,O$Y#s��<<��#$�1!�$ Ɨ1`:j=agJV�"3N�:$�Q�V|���36&d4+6�4|O��a�I8O����Fj�g�<;��܃�ĢoNrx
r&r\0�%�韺}�&ݼ6r��a
���"OT�ȃ�-`���a)�)�ܠ�D��|�8p��.XqO�S.� �EGy��:b���/��X5D^�m`�hW̟X�6	�� �!	���&��Oǌ�uFRm��B��"I)��ňD�� �eŒ	Pƅ�1I7�I(��� |����H0�J$�1̃O���1A�6k	���4��+��)ѭ!�,y`Э�)��T��l�jTz`g؄'�勀�1%/̐�B�V�G��LZtjL��?Q�����S�'���"�)-�*I8q�L�^�R�����?�v���Sg��q$�y��2�i�!2���+Ҥ��d��7��mQ�gc<l��>�ʟ�D�T�m�I�1��k��:,u����I$\���bP�V+ܡ�V�w�P� ӓ:k�f��FY2Qa��� c��[f��!F|1k�-5x2Nۙ%�.-��hO~��$��Mt|(�"�'wI�����$Y=*�RCA�#S��Or0t�%���F����b�/�1ڕ��dQj�o�9X��9�'��'��Ua�#�����nk�c�@�^d�z�L��e��2.@R����O��A�e]�>����c����SЩ���(��A_�� ���
�rD�������䊤+r�3Ll��Q�Zջ�	W�B�L�I:��Q�!EP�p(@Ą�촤�	5[���T9���A=uh��:�-ӋE�b���*ϦW��Q�n_Lx���p*ΤS���.R�:�O�*&O΄��Ag�"DRԨ��x��\�;�4s����i��'>x6$CO:f|A2k.+g,e���'��}�"d�#;hj���
�
�XL�O�x�T9�������>]p��`��U��jJ�������Kg��"=x��O /����X/�xE��O8yc�, t0�:Qc���!���FM�DũZ��-:C�1��3����(D
�*ݧS3Vu0FJ�(��!�_�0��D*���O(I��%Z!l#؄S�E^�[��0$D��آ�2�=�O4�i'�,[Qи���QDv��9�I�6B@̰�>�w��fy���,b!�刺#�
�2_C �#��5@�&Lc�YF�<�IT�1�apVc�,�f�9'��ND�/O���a�U�@����LNjMp���.3/��'���Z��T�]jfC�.!��뉛%!���T�[(Dx@�GcJ�,:ρ+B���! 5;p&p�P�O\h���.A��؃7��|�?i�F )�NL˴��$ ��}Yq` z�:r��:4M�v� I��jK��$ Γ���L� pp�(Mi��hB$�|ӈ���"�p?1��;l� 8r��>e��8e-�3����B�Y8��׮���'Q(��W�OV���;+n�-3���)��$�!��b%��+t6Sǖ�&��ҁ��Hހ��y��	Lր�Bo�q�l�k6��]�H��`U�j�d�&[qXI��O9JuA�I$\O�����C���ye���� L�h"��E�itR9G3P�ZR�i�D�#��Q7a�@(�`��
������2tðU�1��!0���ϭ^��	�!��	��@�=�n�`rd	�!X*#=!D����6|a��لHXƝ�%L/T:�{%�'ڽ*�.ו��s�HX}��i��͋Rmr\�$�'��"��q�1�F�b�>!�ë�4��p{æ;�Oޱ��D�:e�����8g��0(���pt�k�'�1OƴC�Eͨg��8i@�QM4�q�S�;w)�7澸�C�K�]����R';�3"�sg�+~���1�>n���	""�,�$�B�j�	1�V�i���"N��0jʍtS$'?�d0��ZP!v�Ϛp�xy������$h�K�օ��Ë$W�2sp�s�X��ϵ`|s�jJ�|et�؃H��N�]����qԆA�D^�`�n��)Z�E�f�Ce$�����I�Z c&���`Y'71.�(!LʟdOI" Ҷ��?ٲIђ�6���Ȇ�U��L��8M����f�*8lIZ��$�p>YBK9�ưK@��0�����X�'���XG&�<҉$>��F�L0j_0]D��<
�LV�+D�ċFH�5]��L��!>p~�J�ͧ<A�I�p��;4#Lu~��	�����Y ��B��,$;!��Y35��!%��jR���$m�����O��CA� �P��qO���$߇~�6���L)HVx]��O��J�#M�9��1{Q(��bĉ�:%��sV����p?A�Lt1"A���1<T�;肗������Ib��N`�%��VI.��R!h�k�<��M��?�� ���JX�A�n�<��۲�B��fǌ�H�6����B�<6�ҳW�0�f�Q�� ��R|�<a'��:��5���\�
��<��Px�<f
P�7�S ��#��,�FL_N�<�EL��%=��YQn[,� ��u�<�cүb.0q*�]$B��OYt�<YT��Āh 猐5W"�z�)OV�<q�F��v�D�)�j�R�@sbXz�<	C��l��P���u���m^�<Y�X*BS�#� {�4���`�<�.� XR�Xj0��IZ��*E �\�<i���4��]sQ�O�P���V��[�<9�d�4u�<��-�}�ڔ�C	S�<��\L@∊Wǐ�O��=��L�<���U�9�@臞G{&���M}�<A ��[���!��EC��MU�<!���t�~t�D�ֻ	��XƯ�F�<�7BL-5n���&�! !��kA(�C�<A���JVdEb˒ kp$�GkC�<I��/oބ
��ނ,R4cV�A�<���� Qlq���cE�:�A�B�<���@��t�Sd��8���IC%x�<�����$��b�,Ȭw|(!��q�<�� [x{<�'�Q�(��#��m�<��N��O ��������"u��g�<ђ��l��xis�]�V@B�ɘl�<�c�i�Ys��
�Y��y�Gr�<�pˊ�8�|�`�˗�.��=Q���H�<���>�����oK�x�,�GVL�<�o�]��1��]�e&as�
F�<��)��fo��� #�B�^1��B�<��(
Z�Ar�?Q񺔨S��<��G�-/�$��c�7aH���y�<)���&��c�-D<A�c��q�<��kڗc�]sbD��c�|0`��	k�<��ߡPU,���d�te�e�<9Bh���  �D��5�p!s�F�<��Ĥ:�Xxd˂�-�9�P��F�<�+�<X2�-�����2�;"�[�<1	T�@�$��ĒT�n��%��V�<�%D��2�}�BC<(��qH�S�<� �� ^�]��a�%a�k#�\�e"O�e�� \4:,zcF� .1т"O��"��1tY$�ZY��aF�}�<)�Ʌ]�0�x+��|4v!6�Tv�<����[/ h��S�`�d��u�<�T��<�%���X��9Y�A q�<	����{z��*��u?���v�@x�<9�(�^[�ځC
u?�)
p�Uw�<��ŏA:xA{�nԭX%&�G�<�U��) 9!�I[�3���F�C�<sf�:k4�����8(��e��l~�<���C$Q��H!r��rP-[c�H}�<�`�;�����V�
P�f�_v�<IA��b�Lpy&��=^L4a�ufCr�<Ag�U�}�$tN��H7�t�q��V�<Ie�D/����iҋ�py��lR�<��;��5)cFl �H��K�<!�A�:
���/�=.�ᘶ�P�<��a[Iq��+bgζ)j�I�CQ�<IQj@�4�T-�ܴC��7gFJ�<�&T�;3�rì&��M
'��\�<9g&\�8���d��Fn�}	��p�<�ѠӮL�F,Qɒ�3ԬH�`d	p�<��@�$j�H�;|QX��Nf�<���r��1��6�0Mx���d�<Q�� 6���*��ŲI�l���F�<�֧�4�|���jJ$p���S��C�<�"�74�&@`4��;�pA�[�<aG,�a��|�&�ܷ}�����X�<�caҪ���iwiԞ5�"��l�<��^�X7V=� /cǘ�1��f�<a�ǂz920��-�.�ʑi@&~�<���jP~� �K��7����S�<	�M�-Ґ���G
%N4��
]y�<���ڎ)����c�I�nл�N�<�ԣ�Lq��{�Ä�~�{%�A�<1�`�3i ��.�{����Gc�Q<���s �yA����Իcd`���ȓk~J�Z��U�N��c�
\o~���	R�'���0mR$�L<���>�@ܑ	�'��<37A[�(g�H��F�A��p�'5�I�A��?z�,q��ID�d@!��'ڶhxQ��Ly�#M�+*���'ֈke!�"X��^��Y�'�lj���b�R} 4(��lh\�
�'P���) `
 TN��s`��
�'|pq�j�.F%�B��O��p�	�'4�k�#�K���b"O
[�d�'~R�pg�E�k��9�dK�@��4��'�r�q�޻0(���4���'4T��E-_ȾBc)uUZ���'��\�7�J�j%� ����d�d��'�&����"q75�� �&3\D�r�'qd�1*F3P�H���Ǐw~�!�'�AaS \2y( 0V*Ÿp�x�'�̑5��d^.�s5l�R|�C�'��,`e�A�V@:�4ł�X�f$:�'��d�d����|�t���'�.���Ϙ3��m��菱 O.��	�'\�,�"���{�f��bd�D	�'!m��dº�j��N��U���'��L��V0d˶pXCe�O�:��'��ёj�i�6�q2KÌI��� �'��-���MA��a儌?I@Nl���� ��aw-J1�h��K�)CuX1b�"O�`��/ޮ�Ї�)\�m�"Ob����%G�T�ɒ 0C����"O����	�!����0I8���"O�k�̟2��5��m�//(Uh1"OF�D�T�g��i��܆LZ�	E"O@×���` �M�|�$�"O�-�תE-I��ؠG�0[B�8��"O���t�	P�X�l�*E$|��"O��R���=\������C�c� R"O�Rr�B�҄�ٌ7�v�9�"O\YRv⌭:^|��V��=���A"O�H��^�����LHd�*�9r"O\eP���� �^�^��\��"OnT+��19�̤A+Y�t���)�"O��`�ܺD�H�*d
ݽ_�\�c�"O^|��	=Z�x��P���q���R�"O.PZ a�

8���DJI5VE���Q"Oh�Rπ]g��*	�,z��TAU"OF�:��J�Z�V
&�^�A"OhE2�(Wc@�$!���z���"Ov	h��::ʨ@@ F3K��2!"O���iD?J��4.ǩ ��+�"O|2�Dոr1�)eK��>��0�T"O�a�F�� ���w��4�X�z�"O�d:��)X�%k׫7;>N�[�"O�xQ�K՝Q�61�EM
�s$0�%"O֤3�)�7hBF`#���"ԛ�"O��H��()���0	��#0"O�l���H6,�i��·��%P�"O���Dُvf}!嘚u�N���"O�U2Gc��\��%�	 l�e�A"O�k�
Q'\��9Ra��"O\A���D�C��{� ��t<�q"O�q�BCXz������Z,�"O�	i���l��  ��W|}Y "O�ѫ���g���i�j�/,
��ґ"OZ�C�NM�fWH���F�&��Ȳ�"O�`�C�qڵ�"���\6A��"O��`!�8^�L�S��CH� �2�"O�Y�Jؠ]��� ���Q�@ ӧ"O&�C��S'ȹx5�>��D�!�W�/�J쀑ʏ� �l�y.(E�!�`J�8a���S���1L�v!�dJ.w@F8*����&/�E��,��/�!��V>��x��D�6!԰�$A� �!�D Bi�ݻ4�_؝�*��!��Y
�V���	�$���ՈN	d�!�d�)%�ؑ�B� A����!�]I>!�D�OF��cV �$"ζRq ��!�$8]!J��R���Y�	K"�!�dN<r�l����[;���Ys/\<C�!��.o*챔I������ �#!�Ҋ(uN(��GA�*��݂,��=Ǡ��T�.$�0�	$IX�����=Uv*d皹Qu�Aa��a�2�ȓS�\]:�&�S{N՚	^�W�|��M2�[���d�*�:��ߴp������]�JǛ6}&Ų�!2�6��ȓ���"�9��<��lM���|��+np�j�kA-N��5��oM�\S*4�ȓo��8(�*���DP`�I�"g$����`�Li�-�3)$�u`����u��ɇȓhX�!!�d�)T�P��Ĕ5Q9\��S�? Is2� A�|����[-��}Q�"OX�Bi��^�ȂÖ>��=��"OZ�b����Z���a��_�)J�"OX�є�K�� ��V���x�"O�p�@_� |�ړ+Ղ&-c�"O���dI<4-N�+�*ݍ\�*��"O���ď0N�Xj1*�`�^Q2�"OΑ�N����MHDGY�8۶U��"O�l�����;�8)Z���96��Y��"O:��C,��Я���\+�oYj�<���[�|��� ��6D 8��aTh�<�e������E� �~�ڡ�N�<���"pi�D�q��%:��8ڷ/�H�<�H8ar��p����!� g�`�<9��8F��k��$g�"	�À`�<��0z��0��!���E��w�<9a#r���
&T)h���t�<�Sꅵ�&;$f:w)8���s�<�� J�V1&$!� ^<��K�"�m�<� "w�4��K������Ll�<�[.ъEA���)�@X3T�i�<�խM>%�����)OҘ�C�h�<�u�Hx2F�QmK�G��a۰�e�<�S+�{�(���C�}��Q�Ôj�<�+�H� ٗ�N�w��(�G�a�<��ڃB=Ȕ"`�;WjD��][�<�3-�N� kq� %��%��^�<��m�>f��[#�@"dj�0b��@�<v�.=�&��W��3*D��g��R�<����*C-���P���lX�G�K�<I�
�F�J����֘�����BD�<q�#	�s18�&׿A���� ��~�<A� �6������Q8.�P�"�N|�<�Ul̾/�l�ѓh�2hH�P"'�]�<5�V���xx��2x���A�^�<�b�Q=iR ���M�+Hc�Xh�EU]�<i�`ƹfq��ɵ'��N���$�Z�<��k�596�����#r1�l�0��_�<I7Ș�%��Ө�N4�z�g�\�<�"lZ�<��ik��I�4arn�X�<Afޤ��;c#�pb^��[dC䉒�u���k���RC�+�B�Ɍg��4zgj��c6BL��n��%B�	"^"۶oC���%��h@�dO�C�I*Y�"(�b����St���P;�B�	 v#���Q)��XP.Þq�B�ɫ@�0P�Af��pAV�E�PX�B�II$Z1P��B�I�h��Ύs$�C��~�&严�Զ\b��J7k��C��^�H�KE��3������*G�fB�I�!=�i� �JH���2��@�-w�C�I�z�n(I�d�� KWC�%�xC�I %vp��[�o�D�ۓ��W�B�I�eh�����Ou6rɈ�� �rB�	�x�B�R�m?u	|X��K �V)ZB䉠��T�s�XM)X�a�Á�yR@B�ɠX�܉���0&q"�yr�߈FJ�B��P�&I�4��0g �{DN�4d�C�	���	#0�جH��aA&�_�QtC�I6u��X�D�	�rA��K��LC�I{p�A�$E��p�z�x�C�� 
�j ��MK�%E2E2D��
C����Ea�K;dʅ��'��^N�B䉕.)�R&+��j3�U=�B�)� *i�2��&?�6�Δr~�q"O��f*��&0� -�`�x��"OFA9�� �%�BК��(R�%��"OJ4�5k�9Nz����,Y��H:5"OdTX�j]3p���ȡc��x�$�R"O����B[�s��L���X��	`�"O
��@�;qr
�[�@9��X�f"O�a��Ť&춍)©��^���W"Oڌ8D���/���AӔ&�B�"OX�KW�%W|@YEoP�c�����"OXp�UN�8^X�pS�W^���"ONM@$dǶN9D��ƫ�7W���/�!�DUB�XB�
\�\�n��A_�6�!�$�4.���3�b�8�0�D�!z!�䎓Y��<�ǋD>�pi���?_!��'�r�PT��'1���8�- �x�!�$��4���o)��J��q��ճ/9!�[-zV�=b�gJ>�x4i�j��-!��RQ�u��� ,�PZ�
Vi!���*e�Ш#�H=S�"(�*�*]!��c� @Z�+�� �d��@D!�Mq����� ���s�9*!�V�LհU�e%V5�  H����!�Vz"H��ƹ+%n�(S�!�d��w�Փ4N�T| ��E��=|�!�^/C���`Ǵ����[�Ucl�[�'x�*�e @x\����E�p��'��)��LP/l˶�(r��6F�h	��'|�r�l&R�<�:1��>�A�'8^���"ezx8R��!6�zp��'N��(�lE�f��cA�X�����'�.m���� �I� ��^M��h
�'Ċ���c�9��=!A�ȆOZr	��'W��B���G
<�AP��O����'�d�)�$O�TUC��ךJ��m;�'34�A�c�-O���fJ�o� ��'�8���J���u���Q�z~1�'�BY �*��EB�\v��>r\ �@�'j�D۔ř�2�H�1�]�}[��]�H�c�$ψX)t�����ژ��%��tr� �95@<ɷ�_ 	n4��9ô����L�+���3�Fnܘ�D{��'�
�P��I0g.l:qL N��h
�'��8��p�ܬh·��а��']�Ta�.W6~���S$�Z>Fs�Ш�'>Ȱ��*
�i�J��-�05��|���a@��0jIp�Sv�O>�>T��	j��j=
a�gcM�?� �3��	Np���z<!j��O�Ԑ�v'2L@�`L}�<Y�Tr��)�c�+7q���}�<9s��zTvPYEkȤKվ�@5J�w�<Ad��.�b����F���a��u�'say��:_(ؙU��.B{�A��?�'y�0��A�"0�D�#j��/LtI�'�J��LYT���"HX�pw�5��'�ZH7>,��|�%�epA �'Dў"~��C�
i[�=���@�����j�<���].� ݒ��
:��r��<��ѻ?����Ν�t�Ĵq�C�y�<��g��[������P���ᡱDs�<��Oգ� ,�з@C�p�b�Jm�<�3"L�n�V����_�u����D�<w藏)-HF'#^0���*
�<�G��k��A��h +�a�w�<� �� ��6
4�

QS�"O Ȕ���=p�@R��9bP�"O�3� E	mʞ ���9薙�"O>"��;�,z��&#�B}:�"OUKF��3d�ܣ��q#|h�#"O&���[�{g��i�ću!
�J"O ��u!E�%8|2r�R&kbL�"O�	�����r�a�,Y��"On��a.R6#h���?G|���"O��3W&�"���"S�I�H�Hx�`"Ob�8F�P�D�nL�0i�l�vT("O ��B�~�$ ��I��4��'��ɞa$�a� ߇9	 ah4C� I}�B��<J|��ckX��0f�� X�B�I�\'\0'�E;>��H��!��L)<B�I2\���u�'3��1��P( �B�	�t����j�-D�nH�!e_��B�!�µ��O2s88�#�@v/dC�I>o��tsC!�)pV1�&R+=2C�	}��!����@�T�ۣ��Y�B�	����D
Ag�z�H D9�B��+R6�0����������:u�B��&8��0&f�mO�E�$&=4�BB�	�`<F�0u=73��i�fW'pS$B�	�l}4��L-v�X���|�,B�ɋdZ=Q�V55����E.F�r�<C䉜66�c ��LR�����îF��C��t�
p"�0P��5m��-��#<q���?��ƚ8I �DC�n�� Iam8D�����8`�� )��ϋ �����4D� �ƌ�;�F��t� b>���ť2D����ph��	N�<�H��Bc^��y�ôdA�AEH?	�X�傎�y�/�e��y9��Uj*��A�:�?��'�dH��S�2 ��;
N!�'O�|{���^�*�ag�7{v�'Q���!�
�X&�l��H<n�ܭ#�'0�C!! �>=٥f�e� ��'D
��c�-�9�C\�F�.�z�'i�)��*N�V�(r�ɼg��4
�'�0iP� ��
̎���I�83}Y�	�'��h��f�oJ�hA�J=#?Z� �'n���.�p�la�Q��,����'�d�r��l���1#��U��*�'W��(��0d�l(#!�ÀV$���'��)����:<��ga%VT(�;�'��X��
�!wr�i� ŏT��hR�'�&�����%f� Qඏ��_\.�`�'����t�6%q�%��ݸG�\�q�'���"�K/P]�S@N3�|E�'~tٓ�A 7r�B�C�/�)
�.`0�'}(���܊AP���,��Vb(:�'�RRa
E�_�]��&�x���
�'��
��	9Aʔ�����:���'F�T9��,t�8�(���0dLX�'0��*�M�6  ({��؈����
�'����Gj�4�|�5i��pT
�'jL�1�/��t�)�J��/���	�')���D�������K��2x�!K	�'�8A�Oxh�� 0'g(�
	�'��4���\����hVN[�'������@�5�3B@�Zq4��'G�S)] #�z�{c��:!̂e�'e�E��
$E�g�عE^( ���� �|�(�:F�U�Q�(k4�I"OJ@����xKT���n-Q�e��"O�MH%e�
e|Z��(L"e5�"O��f��'#���V��F8���"O(��R�!$@&3d,äMN�yR&"Op��D�O��ɨ��#�t�a"O�Ue��o{��K�k�`L�@�"Oʍ�$C
�U��(�i�"�NUYr"O���!��';^9��iL����"Od	Ѐ'����ѓƭ!���%"O�hq�oC.�"С4�G�B�na�"OBm�d
ʣ2��P%	�W���:u"O�)��ó"ԂIr���;��t�0"O�5���r��Px6����("�"O2���_���
V�V6��D"O�K#H�B�X5���7�܁
�"O�D9QV�q��\�-�2r12p"O�P�)ҬAm�,��끵M*��"ODpX���8x6X��G�"��"OT�J�EE�(��#[�\��E��"Ot�Z3@��M{ ��D�-!xUP"O�L���{�~�2po߮Ou��hQ"O���%�8 ����k�k�@�"O0�Ѳ�5.M��q�k�/
n����Is���)I�D�T���/�+����o	i�!���~�ze*g���r9S.	C�!��3���B� dKv1�@ԃ:�!�9.c����X<`H"!��K{!�D�'D6�hՎT� �tKѤ��k!�D����X��-�-��'� pC!�$W�b2��5��ZJ6qcJ��|:!�$Æ4�ȴ�/�<���΁~5!�$ 0<8��h�<BYU-��w@!�DĻxx4ۣ�I/~\����T=!�V���32�Mv�%�
q�!�D����:�J^�|r���)��V\!򄆆0W "0��4j�;Bu��'Q�zr����h�������4��'���e@�w�x�3iI�~�v�
�'�xAR%�+/�XJB U��2�)
�'v$,��G�J�� \�
:ڡ*�'�:�#��
"������l���ʓo�z x�� �����'3I��5�ȓTr�#�!��JY�Q&ӯ?kf��!u"�3�K?> ]S �-�l��=WT<P5/P2�R��1�^6�
U��m根I�&�V��t!�ڂ�dQ��Q��8�`�pD�a��;.�4!�ȓS �Y���:`� �XD��=�tч�!m<H�鑸?ud�)b	�NI���O�v԰TC@)�XxQ"K�*���g�j��DB�45 �B��S�Z����f����������s�b�7'.�ȓ8?��؇c�;x��Y��H2;h���W���ǉ�9I�h@ք��B�(x����!b2d��:1��^� ���y��,J�lq�pkӥ��$Ņȓb�Xy*��F� �
xx�Ŕ,Âфȓ>�8ay��ע}P(شF�
'Z8��x줻 㑽Y�x6)I�'����|KC�Q&r����7C|֙��.:0P�bH�h��4�pÛ1�ܨ�ȓ2chI	t�������:μ���r��Jqĉ�y!Lu5����8���S�? �,��*\+��!�m��"O �����������p�e��"O�Yi���xF� R�À3�B`;�"O� i�J�q@jX��E�̒�e"O�1Ie �r�� ��d ��I�g"O�51F�@0sQ������Sf�6#�!��ٳ:Ά9S�K2<��x�J5�!�":�	!���F[��q���!� 1s��`aFLEG:�:Uʂ�(�!�dTqѠ,���� ��A%��s�!������P쟍V�ة�TIZ�L�!�ă�p�z�P2ꟈu�|{vM��3M!��҂5$HfO�#xVe鵌ۺ,!� N2���G	�&t�u�U�!�\�v��I�惃*fd0Y֊�%k!�"*hIf��,m�l�"w�!򤇽F�}c!�"`e����G�!!�$%s�<��˽zE�(����P�!�D�ֺ}�H	�m�����
�!�D�	~0����'~u����E�A�!�"��<!��?HA���"=!�$�8_�թE�_�%<�`3�CK�Z!���*f�,�!BGQ�Y�9h^0P!��U���䛐k$T����?4!�C Fc������!Y�34	�8%!�dP�p)t�+���&}�dC��/=!�D$Pv�X!�+Y��X�B	˸CI!�͇�)�'�D��)8Q��[H!�L�	1�L�*[����"Gi�B:!��%#5:0%Ϝ/:܉)iҭs)!��):�p�RL�5q�PZV�(!�ϕG%"\�a�/cbҥ�A� �:�!�O���E����6&Fq��F�(#�!�Ę�xw�lZF��>���E�v!�$K~�hѡ�C�t�F�F�E[!�D�g�l�z�m�%_�xaܴb!�;O�Q%�>j��8@��Y�D�!�$E1V�{�	ܻx����v��&F�!��G'��)�j�
�(�vF 9�!��� c�&���a2[/\ i䮎w�!��M��p!Y���7,NM� �x�!�d�A2�����.T���M���!�D��������?i�ᩅ�٬3z!�B9>Q�k��$o,�9P�A$Yf!�d<m@����B)�pFNؘN!�D^5P��0cP��.=� ��֋YE!���ln��b��!rAjF��.�!��=Z{^����h�"q�ˊ\�!�d�G�
�"��@�E��`_�䫴"OMYbg��h��tG��?�5Z"O�=pSM�0�t�Y�&F�R8�q�"O�,�� Fp.1��>CZ�:&"O��Q�F�} 2�P�b�ޣ�]�!�$]�'Ϥ��`L��K�,&IU��!�$��,�|D�֋��(Dpip��O�k�!��X1bj��+�kN�eB�挲\�!�֋tL���Ȱ~ `�s#�7yu!��S��	��!a������3a!�ȓ{�f�e�,��\xB�S� !�������cGɚN�f�Pf�W!�DT`qda� ��
��!H�eI!��� 6]S������FY�O4!��4?!��+q"КC�����R�!���w^����b�y`P�]I�!�� $����|A Ij_�0��d"O@U� �ne"$`�nϙ�m['"O�p�ř�������*rʙC"O���G�$�`���LU�-����"O��3��le�: �@,�Qa�"O>tA��[���BM3��"O��{�C�.$F�t�f��]͜��A"O�h�&�F f�R�q䉒��ʕ��"O��bgH�^����#O1HT��"Oм#wFؼ% A�$�١I��s"O�L���T�̄�S��#� �"Ol}�j�#�ֱu��dj4Q�D"O�҂$ŷFL��fYAS$бu"O� ���7R�@�@��I,�#v"OlM���H����h��U?���"O<Hr&�ѳ�TZBMF�l#@��E"O(��H�JV^����X�dp���"OJ�{E� ��S�K<+ꀫ�"Op��M�<1��1"PuDl�w"O@�9��ϜLu<�1� �76k�4��"O�܃�U1F[�E#Gb� r�)p�"O�i��#k>d�㎂*��pY�"OH9 Q�O�6��d��d��=�p"O�l#BD�9�� ����d!$��"OhP�^(Q�! �oL�\���
b"O4�� 58 �w�T-;�Duq"O�sk�% 	*8F���Zz�yhu"O�x���Q>��آ��R�-	A"O�>>�{�iQ�t�VQ�SIO�H#!�$��<�F!��Q;��LqP�M>
B!��� >\d%e�'�p1��6(!�$U�?�@���UDFD�$.]�D!��<44ؒ��x1*(B�� �!�[MӰH��K�1%�T*��̕�!�䏡-�X�ŉ�T�� �F�=�!�[=Ro���3��~a|i�JĐR!���%�L��F��bI�=�7C	�fJ!�DW�
��b�V2�I��(2�!�E��PT�g��p�������{�!�$���2=����_��[�b�3�!�c����Ѧ#�F��e�+A�!�dD�����d đ}�hFX
�!򄞈r�|`s��5S�X��QK�;'p!�Ą!��AuJG�i�h�
���SQ!��?��$1F	K*Nx�1�琚vL!�dTF�2�ya�L�s��<	���kG!�$��9pH,9⪅-7�j��;U[!��X�2e�Ǟ.|��!��(N!�
�!����ɦ�Pj���Y6!�$�,8�� F|OD�уK��u�!�d�GmV�'�u8ै�j�Q�!����H<e�̾.R9%K��s!��Ǫ;B�<o�ҭp�Si:���'>TũFj�SlL�2@H�G�P��'�P�(7�Ku3��#�(J�شq�'����_�+c�L��K�.4C��s�'XJMCǡ�
Z���A�> ��'����̵+�R��5"۪T��'j���@3W�ȱ3j(X݉	�'_�` ��!&h ��M>�d��'Ү��u�ˮ.�$�G�͕\�♣�'����2��4^�$S�A��+((�	�'��H�g��_~����# �л	�'��x��B/k$�=���o��%
��� l�Ef��=α�&(G)Kv��3"Ot�V��h�嫓�^�Ek�1�"O��E�Q�y���0�dThrtٶ"O��+b��3{خ�b�!؂px^I
"O��`$��:���11T`0��"O�9�pl��oh�@  �o7��cs"O	(R��R��9%��$^칅"OT�"Q�"ύ�g��E�!Z��:D����ҩI^lH�"!k�0��@�+D�����9!c�#&��7��4BҮ*D�X�P�⠝zU��`1,�{��%D�lP��I����K��
��%g#D�0��Κ!:P�|���Y�A
�X �* D��CF 4#�2q�Ƃ�/�ܑ5+"D��[T�s��R&lޙ_0���a�!D�4�DB�*F�P�(fe�x��e[��,D��
`�(��dp�A��\Z�yc�)D����.�/�(���MF[~u��(D��bD�ůAN�M+�!�>jg��`�+2D�EjXO��9`a��9�1��.D�`۠�օ(�@P���#tDp%D.D��r#�0ZͶ�Y��GD���0D���΅"k�nɱp�Y�|{4	$D��aJȡ$>�]��!�xXp�'D���`cʂ7깢3�ס��}��/D��,l�-z�*#8��2�@�8T;:B�;�"��r��ӂ;`�́
w4B�I�Z��\ٷ˖7ES>T�Wl�	&�@B�	�jhz��'�0bG�L[�F<��C�	?A7��A3A��nΰ(��%?�C�<�@�*��ݔ,���"����C䉠9~�=���Z=�����]	~xhC�I�D a8�	ښ bjd�F�ȶH�RC�
_��GM[ZR���nǹ^6FC�I�O��WHz0U�I3-D,���'�T(jT�L4�*4��ϖU�c�'��@��U��]�ӏJ�E�Z�
�'+�X�퀙y�$�:s�Y8�����'�B�J OǦKPhsl��8r�m�'Ѯ�����P��%�3G��+'Dk
�'	�ːmʵv߄ȡϙ�Yh�� �'I���6eO�h0�5���Oh�19�'t���M�"$\�����ЏNi*0�'(��uj͈h��ͻ�C�i�Z�'c��P��1f$D% 6.��E��'��	[�	ʹ9��Q�U�� [|HH�'b��+�j\+g_�hhP� �"�H�
�'��i4N�w,0�2�n���K�Q�<���	�K��|��m��>�ʬ��E�N�<�j�L���y��X!B&��C��Wb�<!E'J�&�b!��BH.��KC"f�<a%-_�"�3҃��)�`d�wM z�<����c���R�˕:t^*��w�<�c�H�K�dࢀ�2=,V\%\i!�$[44*���*A�Uj�L{�ʜ�:�!�$D�N��3�; D(���ԄU!�d�4>��TG�$&ڥX�(Z�W@!�E�* ���'D[=1���yW-�I�!��W�=l�R6FL�J>�1f���!��{�q�N�C��0�N+:!�$�+B{0Q��f��")� �VB�!���I��[�c4�c��9U!��OJ�0��#M���J�/��
	��yd"O�˷���g�B�1�E��� ��"O� ݋��9�DY�"B�4ǎ��C"O�T[1�_�<=�c�a�-0tRg"O���%OL!q�b��� E�"k��Pa"O*d��&�$m�@<��/aUlYڤ"Ou8�W-���f��e;�}��"O�-Jf�R�la��-�F�95"O��� �ay���F :�hr�"O�(R�GܖX,�;� ��"4���T"OJ���掰_N��`Хb#�l�Q*O"���#*�N\�(U�4��
�'-�26��@�̴hBY�C�h��	�'���!��#d �!h����A���'���"ӣ(�A��	�5�j�@�'�.��&`��(i����;����'�f�8�ꉳ`�n���� -��z�'��L��J	0��0p�I%�6� �'�@9�"��Y6���G�.f%
�'n�a�L�|�|	��T�"�>H��'�ґ��L̙�b��Ū^�cX~Is�'3A;�\�s:�U)��I7	1\
�'0���-eЭ��`\�)�b�I�'eE�m���v� c螊$�Q�'�@`�6E�T�ABFW�D=ܸ0�'���h�M[���P�Ѕ�.L�9	�'7����?w��oB�Y���Z�'b��	���UW�h�U��
��
�'H���'0��D)U�E(��j�'�.��[H��@LI��� ��&�y�+�:G�Ps��(H*&�Ӗ T.�y�bFOjd�bF�����Q0�yR�	5�t�c��?������1�y���?��a'�ΌD��A5�&�y���j2�b���4|������yBa�`j�����_�'fz�R��#�yb��z����e�. �̓���y�27�l�"4nɢ׊���L��yk6���K�h�]��D����?�y�D.o�֥,H��0a�#�y�Cݎ+lB��fۥMֆ�0�R5�yR�	7*�\m��)�?F��ٰdƫ�yb%)}����C #Q*x�'���yB�S�G�,<)G는j��a2�U�y�1qJ���
+[$ r���y�@"Z�^��%^Onֱ�a옃�yB��!�^|��IB�B	�����@.�y�y�1S�@���H�k^9�y҈�]xA˱��!>E�!@����y�#Һlh�d��,S�!���R���3�yr���
*�2oG�	�����.Ќ�y"E�{d�ʡ��UNy�Q���yrIbZR��F��~n�%)i��y���!	]��
��g���d��y�m�N��\Q��_���i��P��y�前Ȭjc��;,>jg���y"F� C���AW�C) ô��Vm���yo
�C_�5��+ĩ������y��S�7�.��E/E ���Y�a�?�y��.A��))@Б��	��y��R=�}�f�U2(N"�pk���y�(P���Q����ԡ"���y�J3Y7�!���ֵ^ʊ� "�*�yh�c���R��ȅM���1��y���E:��S L:A��S`�y"Ep���IFN�@�>��ꅲ�y
� @KW��#0z�i�Aҝ���k2"O�cgC�MW��zTkH'`ޢ0xg"OؘBdiǈ
���`u�I�4�8�"O�k�g�.T� 	��)*���"O U`�J�t���k����"OF�U��#����T%Ls��=(#"O��xEC	3*��T�M'P�2()�"O�����y��I�#f͕]���"O��DoЪ{D�,#3EEo	��(�"Ob̃t��q �cNڂ[BŨ�"O�Ux$�Q��0�!V�G���0"O�� �ƦnhB(��l$��08v"O~a� `V�q��x�A�;Xr1��"OD�)p��G_�Pht�ǣG�tS�"O�M�V�C�MҶe[�KFL��"O��ȅD~�f����l,D���2�FW<<�E�C�r0�fL!D��X�T�����Ɓn��Vj D�x���O/b��T
Fa>V��]rf� D�L 7��)`�ܝ#@)\��qW�!D�p�7�C��e�[;�d���>D��(��Ĭ5];�N�9�,D��F;D�����8�`��4��5RTbq&D��3t��1(9@x(V�N�Y�N�8��%D�T붣K=�,t"5�WH6�
S�%D��A�D��X��@s�BER(�y� $D��ɖL sl����t9(4`#D�8���r�	j�B #=�;�O?D��8t��F��pjgIʈv��)K?D�,�$A#��U�4�	� �xHn7D�|�s���}p*I�d� ߈(;b�2D�\��{-��s���'�"�hrM+D�D	���V
)AF!ՌqI��	�"(D�4��H��B�^)k~<)��>�B�	
z�X�#ӏ��C$�ɢc��C�
]0�"b_>6�P�	�Nf�B�	�Da�aꡦ�	g� !�c�#O�6B�ɳD���S�^�@�0OǔJbC�ɯh|,<x镡b�z��Ǚ' �C�IzH�U �ET�5�:����Y�0��B��l	|�
��ѭqF֝*eە`n�B�7=���6AF�/�΅JQ����C�	�G�\@�f*	0B��uc�U}{\C�	*μx�D�� j��3��!#�6C䉎~��iÂ�24�:�v,� �C�	�\̀�UdF.4�y�dT*�B�I0��DA`[�~0��B�@��	@���X�C��3t��	@/�F[<�+�*D��� aLE������,�P�`�(D����IC�J#�� $�B�H��'D��7� Z��Iic/Ę*�jYjc3D������1Mdiӥ�3g�R���?D��
�&X+ʥ{� �}R��=D�b�)w`kG�V��
2.D�83�,^�JDV #E�:���0a!&D�L����Mf8iRR�C!C`b2E%D��ˣ��M��	c]{u�� $&D��J��d�X��1��+6X�
Q0D�l�+�-q����4`�Y���/D�(�7��
L���%"�r�Q�:D��`���Gpܹ�a]�<�6qI#�6D� ��oQ�s���bǇ�8B�2��o9D�`+g#̐!��u��CO�>:����3D��#�$��*AhvML������7D�� *!9��r�b5Ate' z���"Or8�7��G0��R2f[vR|B�"O<��V�ss��*�e��"�P-�p"O>��q(L<Wa0!1T�J�C�
VLA�<�ը�(�|�2b
�w�No�!�dD6@F]���,E�x�Ä�E�!�U�XJH�:��v+j�y#ڭ�!�D�dm�xB�4/r�T��#�!�dI"<��pq�.ߌB�)��A��!�DNwtdx��� #��=y��d!�[�J��R�	��vΠ�@I�3f�!�$ GJ`/��|_�Ez�G�t�!�P�-����3J�L��e�< �!�d�_��!	Q��<1�A��ƍ�zp!�96�΁"(J���Z�Y!��9/| Y5���eԵ0UD�Tb!�DY�&xL�[��?cs,�WCQ1�!�VN�|�a�1b��a�q�e�!��y�vh3&D<S�����ڦt!�DO�.��{�A!^�Ɋ�'Ga!�D�(�����)^Z$��K�R!��/-�d��͛�@S�Lj���U�!��*pH�P�<{�N��$�B0�!��7߶�US�>�R���,V -F!�$�2/l����)c�"��ыͩ,3!�6w\�؃��L��$�!k�3�!�D��/�z!šƌY�`�C�;�!�D"P
DXW�BmѾ��5�ފ7�!�$�%&BH�����Y�2�;�.�w!�d�78"���GO�l9�'o"C!��-�lyr�E)��(�����!�d��|�V�Ұ�S=̌ÁɩaW!��PJ�m"RF��)\����
B!�d�!R(�{��_��}�!��9r"!��(!�,�� .�f����#�=8�!�d�6�n4��
�ΘQ5lG	3j!�	�Ёc# �a��e���T�!�d����tO�*-~��W��� �!�D�?j�D(	�뉜ªT�VO� �!��mۆ�hԂ\�%H�P�$$� m�!���!����׈^H�z�bdJ/th!���1L�p�B!.T}V&P ��ϟ|8!�䎕d��yQƈ�D^i�w`*
!�dM�'%�!�NY�);����.@/Q�!�H��`A���3h��ch�,�!�d�b:t�b��:���f�(U�!��e��	��1<B��̃w�!�d�?�����O�b�Yp��
;�!�$�(Y��@���"�n0�O/#!�PS�*Z���6��x�D�8gf!�d�VtJ$KBO�7���9�
�I!����U��ڢu�TT�@+��7t�8��J. D����U^�!�wǉ�1Lؘ�ȓLJ�	��D�;	�Ґ����Ԇȓ[]&���onT�H��d�u��J0A衮=~�t�g���@@�ȓ1�tX���_��]��c�Z��)��T =ze�) ]0la$�.�n��ȓ�I3�eM�ohJ���_��p��c���SJ�D��p�Ũ
�R��8qb���[�d���Nv��T�ȓl8lȪ"^bФcPK��p|���ȓZ"İ�̝�$�$���ғSN$�ȓl�a tF�)�>9��D��|���S�? 
"�dˁ[ؐ�Pn��W�0��"O�Ub���Xs�)q�?B��"O�
��:FB�𮄦P�I2�"O0�����jB&҂.��+߼%{a"O`�*T�Jx0 	��?S$�5Xs"O��K�0Qj��E��M��@�"O��2��"]��R�n�> �>�%"Or�9c7:e�msG��&o��y"O�!����!XXj&Кp٣�"O�D#4��.E����f]�4�2�;E"O�t{A/хo�T���^y����"O�ԩ^y/f0ӑ�W�!�"7��b�<AP��A$d�A� �Ws�YQL�t�<)�ƃ
]�PL8 G�x����[q�<�C�rR��gΈ`4�u)��k�<�fO�D>���t���;�]� jUB�<���@�	EJP��49�@E��� �<��c�0F�&y�ej�1[A�Y�B��`�<�ϕ2:���h�/		/J���B�<qN��s��}��m� ��D͂d�<i��X� �:��E~S(-�$"�;�y���yh�ਐ ѹaɒ���y�*Z�7��u�_�%~<�*�']��y2d�����0�ěN���K��y��I5n-1��8��R�O��y�"Q&��tP�d]�8:��g �y2G�l���@(�+q��X��I4�yR�Z�X�!���p�&���y�bRf8� 1��ŝ|Z�5탁�y"�)��mb��X�Q��rT�[��y�8+.��L� 욒a��y���#I�:�H�q|&� �����y�		6E�HA3'��z|�e���y�jV�XR��c��s͞p8"�_?�y�*�_���P_(�XVA�*�P|�'�(�iю��<@"愈�
�n���'9��p�Q�V��U�ą�VY2,��'T~����~$������Ѥ��'����T�
p�p �ƽيp�	�'f�	��'�8b�
d �%A�� ��':v���Aҳ>6�X����xQ�'����͂~���e3f9��"O�X�3fR�vּI�UJŀev�j "O�!��&:J�=���4"O��V��E����v:F��=2�"O��c��<W�V�5��s�H��"O4=��(U�0�)����Lt�$"O�q�dŗ�1�\)�pȚy�"ON���l�l�Nz��ڿz���"O~ �1��53�&-��L$<�A"O��P*��r��î���;r"O`�XB�]�?]���&�ٝ<�ЫC*O�@9��O�P�� �%%��x���'֥����0yx��
O�|J$��'�y�o$�I��b��)���'Oځ���V�����"�(Ե��'O|Q����?B�h�p*5I���s�'�`	��I�6PT�jU��sV�l�'d��FC/7��\XTB��q�h��'݀0�G�GjV�a��f�l���'��i��T�~�)���ؔzP���'�ra��ȧt ��G�Y5�	�'^Z�bmO��E�C gz!��'aT����%���	P=
������� ����b��*�>��'`�+g�04z�"O����$'R�(X"i'4�TDS�"O(XIфW,Y�����.�d"O�d*��0)Tur����#vt�"O�0P[��
���ޜ	k�IK"O�xrcc��P�r��g^v`��Y"O����ϡA� LX���%E^�dB%"O��8b(�M��D�G]��zA"O��^�N�*�Y�!B){�T��"OZ\$�!9&��;C���b�""O�u�ׅ. �6mS�����6�[�"O�4��gQ�����@K�1,�8���"O�؋0Hϭ`�.�������Q"�"O���#��&	��#���%�b�5"O����@��j�l��G2/��	9�"O�|В��9�؋�	Ɩ3��0�6"O<Xr��ٙ0�ZMX�.�d��!�"O>!p�F-'�\â�fh�E
v"O~9��nE Ē�{'��1�BpU"O�u�̙(�8��d�1;����u"O.msw�޺VY�H���T>pv�I�"OT9���=3�(�4c_	1_d��"O���c�'Z��EARj�#�"O��BA�C)n��4��=h�V��"O4��j���,�&*�!?�MY�"Oj��d�D�#����H��4#̍�p"O�s�K�?��%��.����"O.�sԅ�.F.���煈1֭@�"O&����ݏUD���g
�=��p%"O �P`��"f�Y !���-�Hh��"O�8��#n_�pC�B�;�� "Ot����Z4Z�(���� Hԁ"O&|��ӸN��]�4͚.=B�h�"O�(�2�J�0���U'.�*�"O�u�PjE�'��!v&�+[�T��"OjA�!J!8��u#�j^��QF"O�a���j\��� 
N��j�"OjMb���)\Rک�3���@?��c"O Ԙ�NE+e����"//:���"O�í
��Z�����~p����"O��B��]�R�t��z�ݪ�"Ox����
h���.˱JR�ѩ�"On��s`*c}�� "�G�Y>�t��"O���
_���H���970���"O�-��!�&s�v\�$�S���#�"OtpjA�V3��A�-ȏXh�k�"OZ��q���XD*���\]�blg�<��c\Sn]��fٿKp�ᑨ�d�<�6���B{�0@�`�9P'�-�t��a�<A�쑏@?���X�*�ƭ�CD�b�<9ǋ�j�&�����2!v
�����[�<�q�=�pR�¦g#di���V�<��c�1DUЍa�aC�6�ã*�x�<	U�ۊ�N��jV.N󪜫㆘I�<�@��Jm"a0��ʪj�&L���D�<�� �'f����N�t����Kx�<��4Y�����h߭.O��G#�w�<�K�H�v�1b����% 4@�Y�<Y׈өdj�m"b��3�(0Y��OS�<�Z�������|�ȷ�YL�<��.��UcJD��!<L	D��҈�F�<�Q]��H�����)���p�Bm�<d��V��R���?�:��լ�N�<��+�Q�Y��ʙ%XPf�H�<� ��fٽD�Fq*Q9�Ͱ�"O���F#�s����(Ò8TTC"OR�_>X�1�L�i���2�"O��
�-J�%�
�`#*"<s8�@�"O{�p�H�8� ��3Ȉ�����ȓ�D!����nh
=��Z�DІȓ;74�QB♬Z@,�E䔉�lA�ȓ;1j�R��C��2���XC����|�����>�R=��\�Q���ȓLiZ�;�N�1%��; �ٹ~�����7�,�+��I�*1j �7 L����t��m�O	#z�����4R��C剐%����dU�t����1��C䉊j�Lp��h"l�
�FCd��C�.BC:���e�Xp�悋p��C��7^���e�>�e	�aD4;�C�I���S�i��m�8�����JU�C�Ip�9�"ו7�"4+��_9�C�	��,��ba��	XNl�w��#2ʀC�ɮ���K&�@�=�@�:R�OXC�[$d4)�kG6��㨈�9��C�	u� A];!&<3��Э2$�B�I� ��Q�D�$�(�ր�3$��C�IVN�PA�1m^ <�5���a%fB�x-D���	*yR���Ě�Z�4B�	/��yR/��k��q�1d�rB�ɧ��e�QB3V�f�Q��\,~d�B�	�Z�*�YE ��9,��CY�OϴB䉎��Q���$S�@r�9t0�B�I|�t0R(S� ���5��C�	{}�x�ebM�D'�D����C�ɓ%��C`��K�6����S"O�	r2�\�I��\�U�W(\���"O
x*A�O�U��%�0�E7=��t�&"OΔ��_/!�4KE&x�9�"O2d�׬A?��Q��
�v�<�"ORK�LI����Z�NKW��)�w"OF�JB �7╺�oU'n�X�8�"OJ�)%�5wS�yi�B2f���S"O�Dŏ����ڑ�S�|Ǝ��"O�LX�Ne�l�#�A�?
�2�"OF�!.�jN�\���f"O��(7�b�~�B�J6aT��"OF(�ĂËh����@�ʸ"\�4X&"O\dJ�LУs
��5i�uFT�:"O�q��3L�*P˄�<@�f"OD�.��t�F|�ȡl��I��"OL�;Ǉ�)��M9�5��p�w"O���w�֣=�8�k��@�z� �P�"O��zׅm�u�ӧG�0�:��#"O<��q�1ʤ���Ab���G"O�P��V G��+E�sD�<��"ON1* ���h|��rW �T�@)�"O|�rL3U.(Zr$�=e��8p"O��2q���)g��R�(�%{�s"Ov�2i�&g��*sꎮP�A�'"O|5�Q��rv8*��EK��q�"O���6�]�)�>�X�AfT�|0�"O�ӵ�J�)�4IS��.GGj-��"OHj�b��1Sfp��/�/Mڧ"O�9���u�Ġ �*
>(�9�"Oа�(�� X���M�@�e"O2�0J�:o�v�ӡ&��G9h|w"O�����:%���j0��u��	�!"O� ~aC�YjJ�[��O�}ߐ)C"O��H!#Ҭk�Nao�1}O�-+��>D�4A�E�5�\� �H�cw���)>D��Sv�M�8ȩ�0��31,���*7D�Ӓ��J0��:6G����-4D��!J���8�q^N�l�a�g/D�P�`l��c`�hb��3PŠ	�eA!D���1��Ȗ�� B�<zپ��4D��
2F"1�4y҃�Â7ְa�D$D���3H�,�tx���U�P��U($D��:u��R�ꀐ���]+��9��$D��@��/���S�V�Z���e�<D�ࡡƀ��� ��Tv��I!.D���GO-Ngx�&��X�l�b�1D�,�a��E���L�P������*D����)݀�
<�UҺu̴] ӡ*D�<bFI�?~>t9��Q�;����*D�d"ф[*`��[�J8{tri��;D����ĝ�e��a0�ʜr9��6D��:Շ��o�:�) �ıtz���H/D��(���H��8���ޕ7b��iw�,D���� Z��4Sw�sh}K�)?D�t�S� `vr�R���H�1�$�"D��I�,/oY��x�O	�_-Ƥ���!D��	G�V�lz�U`bm�9%�� ��	:D��k�'��%����g�\��˂9D�xT��
���ģ^�č���6D�t(�Bы!�$�7�E�;˔-��3D��8a���P��N��(_P�p�,D�$H��H��d�+0&if<Kr�(D��ٱ=#�� G��p��s� !D�,��ߚ,�@�S�`��t��|0�� D�̫C%M�n���pC�V�Aٲ��*4D��XrL;��Y��@��~�p��0D�PQ	Ѫj�źBa�	.����@.D� C�PY�0"6Ǐ@S�9�4	9D�0 ��,]��Q#-J�9��4D��"���0�u{��@7L�	�J=D�q�
p`u��/j����FM<D���kB/B �ᢀZ�6@�%�;D��"�V<�4�&��_SV��ŉ:D�p�;��P���&k�Fa���=D�xЄ ۻ}N*,Ф!�67E2g7D��;��G�@94�g�M=��s�'D�d��M�VHbwi�3_����3*"D� Y6��H��3A��_� �2�G?D�|A��F>�P�&�8p����fA>D�h�6K�r�����$� 	9�D/D�����%=��!��Y�R*P�g!8D��҂��6�>]�pGԁi(qU�9D������h�v���h�?Q˰�R�<D�`���N�t��W��#Q@�05D���enL��7dT�HGĉ�3D�XG�ʡX� `�,MVQN��!'D�$�AJ���2���>��� D���A���##>��ID���-!
�C��u�j���ժcT(,ЭR3�C�I-�M4)��JtȰtA��n�C�ɯ1�bL�r,A�a���_�/�C�I�*P��V��;�e��'�A�C�	�.)d�1��
(�QSǣT�-nC��"(�,ܱ!䂋KﰡR�$R
P�C��,&�^ё�OQ�j�Q�tgP=z C�ɨ��$@u�N*/L�5��$
�C�)� �H2v��4.������ı_Y� �w"O�%fa-�.�i�*W�!S�T�"O�qHs���_�f��g�X9,��)�S"Of �a����bM\�6Üi@b"Op��s�-$��Q��k�/p�V�#"O8�ReGƴ9�8�6I*��ec$"O��P`���:r��#N��S�����"O�IԬ�4 �[`ҽKm`Đu"Oʉ)��,O@��ɶ�
=8�D0&"O�p��7V�B�H�V3e4��r"Op�I�/R�#"�;��M�	,�,�""Of�Q�hK.I���0�ꀕB*hؒ�"OT�å�/g|�K¯�,%`�b"O�ܢg"փ@��`3O
3^	�\��"O�i�E�0Q�-�nI>,	���@"O$����@�c���Q#ȃ3M����"OzT1�� 2\��R`M�(w7�L��"O�ir�GSy��= �l���p�"O�(8�-�hYZ%�H-$�3�"O��C�ǜ�<,��P��I�"0�YP�"O6ѸХ�,CP���dL̡�<)�"O�I�pa�h�	�@���&"O���/P�r��H
2 ��E�Q�"O��D�8��*��?_��	�"O6�
w" jq�0�o��S�PQ��"O���C��-Oƈ��C�>��b"O����Dd艦��	�)*�"Oh�Kb�"��a��+��oT|�A�"Oİ2K1%j�5�E�^�R8�"O@y��n�{9��I�,�2�ڣ"Oj����r7p��� � "O]xRF�!"�T �&�;~�)5"O� ˶�N�>�<���gh@(�S"OH���� ��&	s���	Uf�a"Oj�Z4kP�A�,u ��� 6*�$"O<j�QAnq@�gL��`S��2D�����z}K��.�J@��5D�T�AƑ�58��G��,��3� D��J��&X�zp�5�:�<��>D��bmnNʼ �O�t���R)D�$a��u��dk����ִ���N�<��CYu~W��E��1(��E�<i*=A�F t�����A�<� ˯-s��1,�"�|�1����<�7�R(�
4�B��&�"����Oy�<i���"S	�m���{�}Y�q�<��'óN�H @$P�T���q�<�5����uS�.��7=4 ��Tk�<�䨓	Ȩ��$iǪg�8�`"d�<a�@�>��n�A��6���y"
��`P����dQ&M����@��yrf�8L-�=�rH۝.I^p���?�y�d\���gC�)A�`k!�8�y2�_� LRYz��°.N��y+Y3: ��e���F}������y"�_�3	��2F��+%Ibl�'�y"�/%���AH�oJ����H��yHC�_�"��l��y&������y���I.�@��!U-���1���y�J<[��L0�O�"���Q`���y�	���x0З��6Y�-��y��)�t�2-�|Ҕ�����y��B��{i��m����p��.�y��U��#q��-\�`c���y
� Pp�ϋ�T�vZ�m��2M�h:�"O���2��
s���FQ�fC�1"O���dm��xW�P�bEeԒU30"O:xb�W�$�B١EH��0�"O�d����L	�ř���i�Yx`"O�5{��7 V��BE�1L�Ո�"OJ���Ɔ�ph�=�'�E?@<yh�"O��� Ӄs�$yU�ˋ3Dဵ"O��6�_�}VF� �ʏ.v ��Y�"O�L
�T�TU �IU�Z@���&"O�8�����Ď�r�	�s��l��"O�{O��K�f����ƙr!.���"O�]s�o�:'�{'(�_�qӶ"O�P�4�P=V�0�JgԈC]�=s1"OX���L�M?v���囤;J�p�U"O�9iSk��y{��0e�n28(�"O�:�i��5���ʧC�g�4��&"OҀ� * k�͞~�` 2"Ot��L�����@�
!2к��"O��;��� V��k���@��T��"Ov��5A�(]�HU�5G!��{V"O`��KZ]2�}SA�[�q��x�"OY7j�)@�zl�.h��3`"Oj�x�L"*��P*�4�xEe"O�}B��	2ʈ�`$�2^�x��P"O`t���J����k0��`��"O�BQǨ6��b4��X&�A{E"O���Ҁ3`��#�7]���"OTh(�#A+c!���B펁&�TL� "O��0�
Bu�iq!" x�F��G"O2%r��>\�.D�t�NQ�ڌ�f"O>A�DW�~8���g��.��]�"O�������*��D�M9�:pv"O�����#$��C�ۚ�&��U"Ox�q��Na\���ʻT@���"OJlxFۊfT9�^��`�P�"O���ūñ~�Y�3�%QWu�&"O�if�y� ����\�=;��"O���J��,{��B�vYj�8s"O��"6��8tc�mx�!ʨy���r"O���D� 5}5l|S1�T;-��)
$"O �VMՐCi�����&t�M1�"O6�A�S�r���c�Z0AZl�)�"O��[fk��鞄ۀ�>dLʼ�B"O�$	3MŚs�ZI�d���0�pʁ"O�(6��(?Qj��TF �%8uK�"OFy��� U�s�T�e{�"O`�6��#A@���C�ݻ~�
x(s"O�xRr��v����E<2J�h�W"O���脸 �̌ ��?#Eܨ�D"O� hd�=Jǐ����,>hpHe"OxD�.�+2I6Ma�Γk*���"O�ȩ�DW�F�P��B j�ɀ"OF����e��u2qX$� @"O��
��k�b��ԫd� ��"OXz�J��&#��`o
�)�F%�"O0<
�Q�F�H`�W�U���"O|@�0&0�^�aC��N��ó"O�Us ��{r>TR&(Y`�@"O�#����n�"B�<~T�a7"OL�Z�MV�m�vB"��I��л�"O��ؑ�r  �Sk��i86���"O�	2��_#~�P�a���  ��"On�#Q&��fּH�Щ�u�x�"O� 0�
4N�Dՙ7��C_�8�"O�q�ɍ/V��u�Ō\"dJ�"O`-y�@��(��px�j�%UMX {"O�U���3Y{N\��jƻ5�@l!�"O�A(#�ߋU�l!�E�{�l`"O4�Eߒ�����dc��!�"O�	T铋��T��$GJ uC�"Oj �I�(��q�p��9m,�D�"O�u+d��9-K�1ː�L&\C���"OB9j�Ǉ2;������BUa���"O�����{%h%��ү9>���"O
lx�#��-A"�HfК1>���1"O�y{�EO
b���"S2،i1S"O�xZB�.9�t)I��Ɗ~�-x�"Otarp�LC�ٻ'���?�D��"O�����ud� ��H���fę�"O�S�@�p�ur��_�`G�d)�"Oj��� 	������+1И��"O����5���Y�iBӠ"O�h��^@��f��AX�3�"Oܨ�KQ�v+�)�%���L��	 �"O�i*�R
' Az��ׅ��AC"O4�@�QD��I7'P1Ur��"O+�V)�B���T��ًpKGc�<	��[�ߦ����G4���DAG�<q"&��!�Q+�6	�Xc֩OD�<�#�Nh��d��x�X��V�<9$�ũx�:H
f���	UԄ8s�]�<1!N�8�� �pBU���d�P
�k�<1�Þ�!���a!!�s�9HG\�<����7�p��H�[�L9�hDX�<C�D֜�띄e4��B�V�<	)J�{�L�
��ԛ>��0uƄ~�<��㌂8, �.�>P������y�<I����i��m1�烄R���cDJN�<��G�F��=��bͷ)���8��B�<��N
�k5r�Qj�*)����@�x�<���ޛ$o4�h�آ2u,�x7h�u�<A`J '/�V���Y p��s�<y�$3�ބX�!<A�.Y���v�<����!G���#"�A>�%���o�<�dHٛ,@ԹAE�$? �s��S�<���15��p��]h�^���j�<�söF�| �6CV�A;�p�A}�<	�bH2<�ܒ�Ɛ!P@�I���b�<�k�O���@o�2/+&Ts6Oa�If8�0(���'`2E����4F�*�R;D��A��U�1[�͛��
PJ�
9D����#\�RM�ɃBת6�lZP*)��hO�Ӎ`niA꜒�l̀1�ڧ�nB�%�A����O0di:�[���%=wў���HO�,9���R �պc$Q�ƚ��!�$�0�n�XL
Fx�<Z@`^� �!�D�g�`Ч�<`�\��ѝo��{b�ڌJC���A�Q�@�y���!򤏾y���
D� �JGj�OjOH�I}�O֜��r��' � jh"O,	QgDL{q@��m�V벍�����?����O��� 7S����O5�̸�"O0a	�@H��V��0J~Θ`�6�d��(O�'��<2%b��g��L2D�/q�(]���� kF�f5�Y0��q��Fz��'��`��K�>$�� .A�4�t���'�Н��AI�g ���$ņ"cj�c�'�
� ��CG&���F�ِ�J� ��jd�'�qOd����J��|6���&�3T"O��q�	I7 �	d�� r�U��'�;���9*�r���0P������)=�$B�2u���Ж�ۖD�Ii
�Y
���5}��'��x�O�r������'&���ち6��a%Ï�ݶ��'�ʁ��	y}�ڡo����'��'�7�0§���C�{�	�J@r:h��$�#341O��{��?y���7Qve�L��UIfӎ8���A�F]��l,�T�P-v�<0
��
4� ��*�a$�فe����DC�q$���k$9��$ɆH� ؑ0�O*P' ��vls�'$�"}��G��y�'�F=R���p��Ա��B�I%tNсWh�.J�aZ!�W#w�VB��7|�9a2	��h̬�� bUL|����S�<1�g̑f��=pC䕯��zC�F�Ĵ��鉹�6����7J:�3G��}��I��HO�m�-�3��&Dç?� b���x�<ib�_<
T��;D��Y6����_m}�Mo�R6\�i>c�ޡU�dH�U��3���HS�!$�L���D�D`b�
��h�ƃ�K�<I��ӝ!B2};Tb[Pv�H�V+M�'�?!0��&��Y�Bk�G�`��!k?��l��0�S��P3<�y3I@tO!�B�I�q��'��fO�1�W�ɦ^�lB�	�52���͞"����� C�ɽ���]2u?�]�U��3��C��'�|+�X	T�*�K0�D�=~�C�'![��H�$r�y���B=�C�I	�fH! l6q��[㌎1n��C�	1kU$�4�bd�UA�4O��C�IL�8�쀩����6��bVB��П�z�@[';�N�˃�T�myb=���$D��5�4FMJD��'�Y���@G�!D�ȑ0I����xUC~�2��/?D��x�/#x6 ���F(
	�7.�>�޴]L�O�>yB�O�U�<�G��?N��k*D�X�W�E5%l8Y��G�*Qzvy�d�&�O��	>a����L�pۆ	�偕:<��B�	צ��fN:g�tX�&��$�Bt�Y}��'�F�(@�H'4o�{=��r"OL�"d �	�������A8%���i�L��	�	J6|�n� W�0TQ��R�U����6n��6��x�k}BiX"R�yr���z0��A#�y"�^0��-��C~l���b$��X�hʓ~��)�'4"U�b>��Q�]�b��XC��>W�r�X�5\O7�#��*l(Lsu
�(u���'D$m(X�@��	%A�����kI�f-��s��@1Z�c�h�O66�/ҧE���W?& ���K�,�xi͓��?y��	{��("D!g0D�����zy�HH`��H����H�˳��"����d��s}�'����*8HxQ�)Kt#P�2C�)��<��M;9�i��"C�`Mke�X�<�g�P�P��09�]��@Z�K�F݄�2��`'�+��1p�né:!DB�FZE��"�$7�=@w*��d0�ɞ��ID~J~�'�6e:�
�1}R�Գ�h�&s1v5ش�hO?7� �p���)$���������,dG�	}~��'N~�:�'�	�(-���Ź4̌�J
�'���ӖG�8<q�����-�M�
�'����b�St�$�3���~�@	�'��S`�̥3��\����
�9	�'@�i��WV7���b@�35��'���C�@�+��	�:������ Xؘ��G�	���٤ʀc"�Z"O9�4j�#��!X
ǳQ����p�O������́W|n$����rŢ��������?��xs�H��}��8%,ï�!�dG�;�)�@"�%o�`(��*F�!��h	�<����{c��KDMc�!�D�N̺YW��;#Q�ʓ)�u�J�l�_����"N�(Gf����/(����0�y��wɨH��)ޫ&��t������'9ў�(��6i=s���#݅k��ە"O<P�2H���h�câ	�,(�"O�y���4a���b��)���#b"O���֙6�9�g)�OĔ��v�i�𤍏=*` �����X��@
X!��Q���b$�ܘ�\�g�=K!��ً)��8�*�.6��L�1��Ą�t�ؽ��ȝ�:Y�1f�2ti@C�	�(t�Z�"�5��ԃ^�hmDz��ꒊه2���f�O(2ޘ	���1D�P;P�Ҙ2��))Ӥ�_\�M�C�Of��hO�����g�(�
5�'�X=����'��I4%J����ץB���[w눗a&C�ɦD���9e�\�_z�u����>r�\#<�r�'�?��PC��h�@a��Բ$3��!�@4D���J��%�� E�ބ<�����O��=���HOfM5��RM��8��UJ�
�"O.�pZ(�ђnB��9�w�*+!�dV??�䠠�ߛe�Ba��(P9a|R�|��6P��W�L�P*S'�9�'E�{r�5$�^e����7.�B��R����x�'��0Ń�s�-�1HҀ�jء�'�\�6 �&/�B��$�I�I�'0��� _�|ͻV�Ρ�P�
�'ߚi���g���y���b���O�����$8>���딶E� �P�ާlTa{�R����:ǰ�����4����b��ai3D�x0�J 2O���H�/X\�R��-��hO�OBՠ!���zA�Dm&4�B�	?*�Т�_p�.m��d*KA�B�I�ItE��˺ \F�˕n�B��72��=`���{xe��h�&J�C�	$U ����F ��csI%I&���z?IJ>"`�5.�\�;6��.v�܀1�s�<����F9�3T�J)C�8��Hl�d"�S�'8dpؔB[�jHL��
5b�܅�xa��h妙5D=��)")\0M2�Ņ�RF�kFAؾW*L����H�ȓi��U`�K(x^T�a��$%A��s�m��WC�}*g��+
$фȓ@	b5�g��d�Ԝ�E!�]D��	����Ҁ	E���I��h�ԇ���Xs���`d��T�L�j�̭�ȓ7WD��a �;+�r�Cn�z�:��ȓN�J��"���A& y�(���r�d�Ia �,	wƩ)�ܾZ�d���y��᳃živ��9v�
�O)�Մ�ZdV�	��@1��L31M�8� %�ȓT5�ph�O�0~Z��D�TR'�)�ȓI��1�	`��C&ͬh��|��As�d��
͵Vf�x
S�ނi� h����SÅ�-P���v��3l�� �ȓU��s#a�'VI�kZQ���T"OƑb#��0<W&�0�%E;K����"On4��h��$�@C������!"O� �����/gjv��e$C�Zp��"O^�1�o^:d|��B��r�x�Yf"O^�[�+3�ՊЮ����c�"O���ff�4{�(�1�S<���"OF��#Ѧ8�~�@ O�f J�b"O4�(�I/n :���7C��D��"O�ȃ�pN�	r�L�8,�IPU"OJ��O�%ĜHR��۵k�����"O)�4l�5Q�"�S L��b��4{�"O�]����L@������u=�Y�""O�U�Η�2�f�@49'T� t"O��s��F��i���1���V"OhT�p̜>"�9����%�l��"O�h�ʞ&I
,`��ҁ/ൡ�"Ob���,]�E%0�%�V5�d�D"O�I���E� �!�;~��pS�"O�h��b���|���}����"O���#N>���(��W�
�R"O�h�a��_����1�U ��)��"O09�p�'F�ܸ�甐L9X�e"O��Aҋ�>�΄��ȶC&l��"O )���Gf
�g�ȽOp���"O�����ۺ�ܜB�ő�ir�%��"O�0�cM����cn�52,��q"Ol��$��Skl��V�Y��r6"O*`8�*?]Nd$�A��p��"O�����.���6�1�><9"O isuD׼G��r��!�J0�"OR ��m8�F��@�Үk�$��"OJ�����,?d~@lōEJ���"Of�9�윇Q�p-�!��=(�DE[�"OfX2�i̚�-���	��x@"O�@�7oϸ~ޜ��h˱J�dqJT"OtY�ǓO F,�T�����p�"O�0{F��+�He�m�X�8�	�"O����'�6N �%��˓�w�P30"O�����A#B��5��& �&e!t"O@
�GQRL���/	�n��t��"OB�k�hN�:rF��m�:r���ٲ"O�h�`��9���� b�vTH�"O�d���훷K�F��a��"ON�I3�ؠ��� p���� "O�Q��\�}7*�S�M�+����"O�]Yl	:d\=ڱ��8���U"O���L�U�zwnE�2v���"O6!�b�.#6��ZU�Q
p6P�"O�qP�Hƪ#,����F�w�Bm��"O�pi��Y,-��P���}� L�v���<�!I�=-�N�����%����$Qp�<y��b���y���J(�[��Jm쓷hO�O}�`�U�䊣u� Br6era�4D��1�q`���#$@ p�j�O&�D�r���OM\l(�b�5-Pݫ@��9Ԫ ��'
XLPBD4��<����:������+<O.|�wj+{��� S,@V�YSf�'|qOU�'�� �P���A	u���H&"OV	����
�Y�b�9۰
�9O���$M 7�ȹ���ݿQ�,�jTMF�?�!�$Ģq��Y�� ިB�l� dL��ly!�D#ER�Ȣ6��3<�N´L\�x@!�Ě�R��&�"{�у˅�?!�Ӵa��LZ��( 
��J�!�N�}@�Ě�K�\�e:�	Ȫ�!�$�dd|�Q@��h�@�
.�O ���?� �����B�2��p��΂��8�*��'��qmZ`e�}u*�1$��BE��~Px�O�=�}�u�^�a/ ��芚u+P�2���H�<	C1<���� %ד��b��O�<���O�R��XY�N0F�0q�FH<qL�)3:�8�"�+�y"?J��HʣQ�h$����'�̝����B�V9h5� 6X���3�'1O���|B��DI 	T�|:eF1N�h��ÄB��p=��}��!4Xf��K&K����`��%@��Dx��b��'2(�O�,`�JX�l�p���GD��IT"O��f�1�T�e�Md�HV"O�I��>:JRI�#��95:�Q��o���)���h�B4�=M����ϯ'�!�d��YY(]���Z�#<�(�
����'m����Zz��G�\#6�R �f.�|�x�@��M���7�@�B�K?��Of�ȋ���
;�]�a؏�,�E�ͅ�Q��E{*�����L$�,�1������#"O�X�P.M,=��$ΜT�����' 1O��d�}����-"+$�QrC�6 !�ėv�̕�4��QL(�	��x� c�8I�ҎC1W��3�]�vX�m{�'5�܈��ʊfT�ۧ�V(t��1q�':�6�)ڧ|� ����9���[2.�@�\F|r��g�N)QF��a��|w�ʎf�ĒO����E!K L+'m��il&YJ'n�j5!��I�^Y��$&�W��E�cq�	�'.�����
Ih���/e��Q��hORY0G��J�
�X��FB��$X"OX(�0��lҌZ%jѠ/Y��XX��l�b��(�r��3�����BќwT��ӧ"O&t�ĉ*H>�!{�ѯx9��՟|��Q��F{ʟt�Q�n�n�  K��x44�9��'��>V7��CŀJ�4m��A�.�B�ɲ�x�qBҸ)L �J��D�C�t�����EK�.K���eg/О��d��$ٳJPI�8K��M�����1b#D�l�b�_A6�X��E0'\f�C=�Ѩ�<,�sa�mj�"��fH1��O��I]�D<�&T�u�p,�,.�D�Y5��k������"v��;'X(��'����n�A�����6��Ej6�A�	�)���`!
��?��'&^|2�`2��Y4�JY���<��D!�OΡ��`�\v=3��)t^�¡�I�MJ?�8������р�o��ٓB.D�$9�Hެ~��؁�CE�w�̘�$2��hO�-D\�$��2� г���U���>��`.�'s�������}f�-�'R��z���`�@�#��0J���{%�Q�%.:��I7R��?�'�O�|R%0!{�Ģ&���,H�q��'��IL~RMP�E�X���Ǔ�8 r"[
�䓸hO�2�D/8�%�#��J�m�6���'����)�Ӧx�>�5B �w)�X  �΋ra&lr��.��"~���uR�`3t�&r�q��˿k��C䉣�؀#��H<A�[ԠI
o��C�ɾ���S��eN��ۗ��˓�0?���� ��u�|f���/�qyB�'A�ɓI1z!"�C�L�|�2�e?C��e����Ѡ�>}|4k�cE:l�B��%���D@�(d���%��Us��PG{J~b��r?Z<�C$ݤ]��m�q�_`�<I�O�_��
6BƤ$~4Ȓ�D�<��#M�i3�F�U����Vi}��'��DGj���:A���1�$Qu�\���8O,c�� ��#���5��Yp���v"!�V��
1��'+�'$�}�Q��t�h(wM0���p�'��O�9�4���떻"�&5bo�f�V����0�'�V�Opq�l��k� a�b�>~�.�KE�'-��I�k�*1Cu��U�^�I��,�B�	I9��ñbш10t�0�)` ���>���܀@ؘ %�>74�pc���=�0>yq�8?�sb�6Q66���k�L�\�03I�u�<�ԃ�Qo�Z�9k����"!�[�'%��E�T+(#w��Ц�h�L��Ӡ���y"e��&_��	FYׂ} ��*�yB�D�������G�]��K!U1�y���gݐ����
\�p�����y�'8c�t��5�1U���EP5�y�ޓ�}ye�βMi.h��y�dR.]���E'�0��A@7�y�M�n�f�8&�N�D�)��$���yR�ۈR�Neaeb��pU�-�D���y"�90�
Y �N�8XF1P�����y��Yf8�
�9A.��� M�y�#υU,,��V��6�H��h�!�yҫі0�Z�9A`�-��,��G��yB�]<&�
A@V�+�l�e#�8�y�F�4t��SwM7y�<�E��y���|`qA�Ԕvm���T�ӹ�y�ާ���l��k�Ѕ���V�y"��t�d��O�-]M�5�R�*�y)A�y�b��7�?s�����V��y�a�Y�
t��"�.�j�)�B�1�y�Ğ�!�\��&����l�Ad��y2��79���.M�^f\���ݎ�y��͒�z�Pć��Kb�(�Q��yB�sB�%�teĹJ��� ��ʽ��IPX�x�P�X��乺2�D�
d;6�#D��u�8I���iB��
=y��-D�|�wl�i��Y�E�ۧS��yjs	̧T��7�)�矈j׆#,T��Q��7��0&-4���4��C�4��-���i��J[A?q�'n�YY  ;M��k��8���r���4��:�`H�9eH�n�	q�C�I?��p�pnѦ& h
TȈ2y�B�I�;��%�oK^��a)�`��Z9�B�	�cK,<��d�1�ډC�L��7�B䉭!����R�~Uh̹���7�nB�ɁvIj��� Q0O�*h��눬uh��ƓYev�Q��!2J���(CV��ȓ'=��*Rˇ)������P��ć�U����ď�zh|[s"Z�Yd�p�ȓ$[��`�C@&'����B����ȓIu��X�n����uSu�L�!`�0�ȓ1 .���ě�&U۰L��Y�ȄȓD�b�[�,I�����W*%��ȓ^Qj��C��F^r���
w6>�ȓla,�#¥��l���s��VZ<f�ȓ��ۂk�>��5��g��l���ȓ2)̀����dT�aʆ,��ȓM����B�@�RF���7G �����w"8���7H$���A�:��ȓD��<�K�"j	�1鏸DL����X��O�%)B�v�&1~y�ȓMRu�r�*:���ݳEi�E��a�`�P��a�dt��M�dގ���V�&=��l[�+S~ �b��=C�Ұ�ȓ �d���ϡD>��j98���S�? D,�7�K���@Yu����"O�x��ϒe ���`�*=�X@@�"Ox9ˢz������&X�4:"O"| 
`8Za*u���$"O<�� NH,�|57"�+�bdS�"O(��I�X�����.Z�gTth�V"O�����'��C�-rK4�8�"O���@Q��>��0↛|��i	�"O<�Aԧ�k��dSt�D����"O�,��FC� ����q�ҋi��qc"O��h`�I4q���2B�F>�1{�'��4[�k��'����m�e̐�r�'���w _ 2t��S�U�W'̔��'���ҴnZ�/�x�Ã�ŦS��p
�'���v,Ӥ.�d�!nH6Lh�@�	�'�lE�2.^���` O�rg
���'T�l�lŰV R�jK�l�����'�����/0\�j�Ń�{�L��'�ʔcU*>�$�{$��+�,	�'�~e� ���f�p��A���0��'���"7�'E� 
ĮI1�ڈ�	�'X�	s���f�� 4�ݢ��l��`7��&��E��{©O )��$:����Ok�B��N4�y��F �Ny(�-@=G�n�B,�y���?ɒ 8Si�:Ԣݚ���y2+M?M|<@�e�2b��hE��y�4��@a������ 2�yR@�=�b�@���$S���ybQ�8��Q��S*���h��y� G�f������:Ag�����y�ܠa�n�ö��V3"��a)���yүV�2��yٕ�L�VHQ�+�+�y��&%���K�9^�U0� 9�y�سh�Yy򣃲?�(�a ��yr���r�&��Q��/�(�raF�y� P�*i|%�	�%�&��v�
�y��
.G�Ф"�,�`��5�P��y��ʘ�b���<Hؐ����|�C��+6頥`�^!&0�TJF�\�"C�I	(㐹�P���k�@��=M(C�I*~��4f�G�k���g�-a� C�	�W��A+NI!}r�#7��nA8C�ɞ`g��[ۥ]��}��O&8?��K�A����S�O^(00������.:j0(R�"OXL$�?�
= aa�pVȁyAŅD��B�!妄+�*����@+~ �^x8XYCE!da2��2/�Xܘ�P&��\��}_� 1I
��q��'�ll�lѮA��!��L/I18��$��f�b%*7O�:Va~�O ��:$�|���K���#C|��2�'.����
���!�Ì�v5��X�ODD�Ŧ�j��1��z>9�g�5}P !'%����!�1D�T���of�5f�/b�~��w���j�����7	��L�9���%>�yҷ�r�	#_d����P�9/za�叞2�"�� ����hghˀY�T{��]b\���	�w�� �E��5�<��s���"�i&���M�k�'���s�g�,ߨP[iƟo�VA�7*K$9�H� /��E�l8��'K~��IR�#(�$��<����G�8���C�I�>�1D�8��	�Ϟ�M�\#*C�D���*�	0U � b�I � y��Ա0�!���p�b$��k *&��e�'��A!��Ɠ;��aЂ<\(X���"=_ʓ�r��rl��o�b鱰���G������v���9w\n��+0E�$� 5B**�ޘc�e� ;��!TK�Q&L����I�\.�&M(���堅�S�����[VDy�+юY>��5���wy2�K&ͅ�d�����^���k��<����/\¬�W�){~9�>�Sꁟ\I�
�L�6n�l9��ߡ��3� t<zfC�ptkP×�M��d�Dӹ;[����9�'1P<t��.�g#�h#@@}�~T0SC{����
2
 ���E�O>����9�|��w�A82&�QF�ٓxR���l)��'�4�|�'�(2�B��)��;E��)��������.���b�O3_����h�8�u��ɯVu�p�u��H=��n��[���z'̶_�����ΔC�'�J)��n%^����G��"��̃�gn(=�tIF�N'�uP��ª0�Q� X��S!M�pL���ǟ���'�U�,����-�Vd��9�I>݈%3BB	*d����԰䧟n ¦�H�'N�	�o������$���ȋj��o���}��S<����K'�@)��O&T45��(��̸�I�P���}��'&XB�Ɣ7�4�	��ʱ+�ԫ�bD�SbXeۇ^�8�#�3�g~����NL1�l��@��f��E�� 0HdY
&
ωc��D�q���3�{�F��0`�W5!A91`M�.$T�`���=?�vIC�d��p�:`�I��p(���g���&��g?���O�v��Y����m4�b���I6�%��e zxҝ�&�I	��d�Im�)�n�&W��q7�G�����@� ��d#�N�LS��t���j�(���Q:3�)�݂�M�w���{_)rf �5#��c 
Ď{נ�|��X�P��N*I���7�
�~��݂��<⨘�D�yw����S��y�i
��x�7��B���`�[����3�
��U��{�˟���먟��GxGM�El��U�$P�#���*p��V
_��cB�Ż�x��g͖Dl���Oڑ@fk̖>f�:+S���E"��
J�h��&�4`�6}kA��$�"?IT��8�����-n �<h熇<
X&,��#@>ش���wjr܋�%�b?���i�c�^��O�r(ks�D?h�`#*]}�ٍ�D���2�O���O��	؄&��I����g��h�� ��4 �ތ�0~���q@���<�'I���㷇C�$�9+E!y��ƇC侘�F+�N{�$�+M6<*�{J|�UDG�8;�yB���Z�v9I��B�A�-��%�6`�	�&(>�K$�P0/_z��	�9V
���,�
�Ek&0m��=�R��D�b�XAk�Ԋ�Ɍ+7�D�E���i�:N�N�� X����'\lDz���"���b��to�-(��F*�A@�ۭu�d�	/2()R�C�q���T�6Ǡm��L�d�n�Kqi>D��
3lم4�i�5Gǚ0�&-k�f�X�`_�X{h�ic������O����c�,�DmZ����0Df5@'K�n3�}"�ˢj9 �����A!ٱ'�Ə}�Uҍ��
`��/��ɁĆ��;8�P1D&N�^�G{�<nu.�Q4�NN�(�N�3kٸi��L�GL �>�Ľ�ȓ�H*� ��R^쉄�P
~��y�2
:| e`E�~���\�7m�S\���
��q���r�΁���UJ¤�f��Gar��
�b�@c[:EaJ%Q$��wd� o֑
1��CDF��F�� ��h�P�O`N-AK�C�]?8G�]��HT76Ql�Rp"�Z&�C�*�52���"ER��V	ܩG =��٢+�i2��h�΁�!Dp>1"�b�!BqO�0j�lH�"  i!o�C�v��g�'� ��]<wS+��H}̬�e�H9h@��E�i<��L�uS�����T��Pp�c��Z��-A��G!@�#;a��I� �F��2;"B׎/G�Dk����	p�S��E�5j|�S�W�&	����,�p�<�WN�B{:����Ŧ�S�%� ���ѓ�NY���+��Z��Y0O�=��|�}�;=�a�Fa;~�ؑ*!G��?�|��s�fm c�\�)H��G҆
�j�#7�V7�܅�$Qnu<]ȐJ��|3Mܺ/D㞜ಫ��]���b���HFE�j;�OU��j��R�BP�u%�dO �CgI�L-�|h� q���y�Dб>|�\�T̆�p=���E�Ne�|�4�3W�jzfDR�'Έ�pr��7������2g���8�,H'�ԹH�Pޤ��D��O߲�c�(�y@q]��@2��k>��'����$8�EH&Qĵ��#�8p�!@�Ls_��>�;� ��A̅o ;B��3Y���zU�E�rJ�2�a �̄�ͪweY+��AA��R��D( ��K6�J�>AR��$D�)O�8�Z�oCu<�� �9lO�}�"�;�)��))x�qr�m�t<h ʕ����&�P�&�C�(P�'�'D�8l�M_=[3�3�6�I�s�Լ�e *�M�-�4|�`�(GȌ�[����(|(ډI���Z����
��y⫃>>�������5]�X3�hV([�.؛[��s榚/x��	S�+U.Z�ᱏ�4jvޕJ�iL2K Z��d뒢�4m)�h9D��[�-� �ŁeCW�N�X�F�T�@��<���]1~��dKŐlsD�]66�p��֕g����u�ײP�,�JT�SDMa{2J$V�>X
�I�)ɦ���D�<.僣�9`��!A��F.+F�p@S==����t�,a��]Cx��ަ
z�b����iB/��U� D�	Tn=�5.O/~�>���Oތ`��L%�E��P���s�\O�<�ō�6�{�E�R�4i��_�R���CиBy.�8��D�J����EM���O+�� 8�piU�z����+�/%�P���"O��r�ń�`S  �׫ͽ�fp�h�t^@�3Fł x���#p��X����aV.�h��/����Ԫ��*���V-bӢ�e�Z��X�?A��ݷl,Q��H�%(yZ( �M!a�����pu�g��"=���	 a����Q+�	�Ĉ,����p�A+#H����(8�����I�be�@Հ!@u�
T\�0
��`�� "����V@̓"���j���j�)��)ك$�E³�U����DM�I���d�Lr���`C�AV����������I�U��<��Lc�P8V�-��l
�M2z{��!>Y�"|�'q��T,�'E�(Y���3Z���.�~�	�?I��X��V� zr�Ef]^��t�Q�DQ����K5Hb�y���H���h4�	�$Z�U:���-a:İy`��
x"���vm?=	�鉼b�D��폜���� �8EcB�FKl����̣@T">�4$��iNj�|�v��A�]���;#�X��H�j�&�p�Ȗ�k� �Ј�i�9Zv\������>�D�&\�3�1O@�6$<<O�,���da�T��+T�)U6`�'O d��qVf�<���\����	�5���WgŐ4�(@ ��(�!�D���܀�ԩ�=ZA�LR&h60��*�O������5|O.�`4o���B�7bP�;!�'���˱-��V�JL͓6�<�h��X;K� H����Z�d��\`Lh�F�(���`�͑�u�>IS���B�t�9���ˌP��SPdݩo �]��"аd�!��A	Yp��Ap�`Rt��_�L�!�F�i���ƀ`Z� �Ήh�!�DY� �����.�٩�S�9a!�DP�rW@�:�L�Xp ���g��GX!��T$��|Ym�$I*�c �O�INAF{���'�bUkR'FL@a�r _�z��|�	�'�����Ϸe5�Q�R��M��0�'a�牴f?��%GO1IE�@�����p>yJ<i�C�<�\�HQk��^ӤX�C�NI�<I��ٹn�K �@"7�L��i�E�'�ў�'.�V�B %-m\���mϽ�!���1���I�@�vg��9C� ��E{���' RD���v��y�R�Y���[�'< �r��v�r)!s ��Y8���'�a�ٴ=��Ҭ�=q*�Eb4�p>�H<�rhPh�C��^U
a�!�Sg�<�Q_�f嚠{��\%4*CCV�<9��/z�hq�p�F~�Ұ��$(D��A� #s1�  �@ �dH���6�%D�����6�R�P�@�W����i6D��� *�%
����
�Q>`��F�3D���BѪ ���Q��)�Hp�/D��1�[�D�����h�O&8��m>D�(�6�@�\�J��j�9?{lx�t�(D��V$�<>��*"a̺}0�cg�0D� �5l�����1�,� ,]��o;D���P��xM�ԊȪ2J�Ѷ;D��BjRxT:M!F��A��dD,D�D��JGK�`�Ǥ5ުUR�-D��1��\,�����I�& ��Cn,D��b�,6k��\2q���FWny���-D���ѣ���>��Xq�Te9�l�8�y�aO*u �T��GK+~���F��yK<#��R����R�0�l�:�y�F�=j�$��zN����)]��y���1$��h#�j[=rK��%�ŕ�y��4&&mk`U jt$���E��y��:�R=@6f�l�Ν�th&�yrjL|(&�Y6�vh�����˞�yA,,��m(����ӭĈ�y2����E3+483f
,/!��6mV$�2�L�r8.YO���'u� *t�<=;�8�$�M1��
��� ��)k��Ӛ�+¬��Jt.�4"O��A��Q�#g��K��Ȅ@dZ��"O �`a��z��ⳋ 4l�D"O���NR"km�A�"��Z�Ę�"OB�U5���$�$xN��"O`P�j�J�Gm
�M���@�"O�]ke�B0Z�� E�
 �dJ"O6`d�_;M
��t�L�!��"O���]�Mi7i�X�c�߽�!��Æ�֭yb�̊c�`|i�o�?t�!�D	����+B=9`� `��)�!��>~\p�˖�0R����M�!��U�m��x��'B��lڲ���v�!�d
%CiqRX:�(\�� ��@!!��H>_e������.S��T��J٧S�!���7#d3Θ8A�\��P��!�!�΂YF p��@P!B�1�Bf��!�D�
dF�شg��':��;TE��g�!�d��	G���7&�)�e��o!��,WHT���	&��03p!��,q;�=�@��W x
�$��!�ĉ/p��
r*�Z������@�!�D+�4c�̅4f���A�!�DV�^/D���,[q�>�Ac!-2}!�ĕE�x9��Ҷ#��|�B�-jG!���B|h��/]x�
��a�c!�$��Q�
a�7�͙�|�[�`Y5G�!�Ď�;]��1A��N5�ċ��N�!�D��3�,%���2��e�&���!򄏶=%�#b�GCe  8��W�!�dP�
9���hD�t���Rj�!�d��0�I8�`ƅ�$51���f!�DL�i���@B�ۼW��a��N�!�d�"	�t���M2U[�]8�QJ�!���&2��(�����N[ �@Vb٬s�!��И�C�@ř7@Hx fk	�|!�DR�r#`��զڌ[4ҽ UɝPZ!�U<$Q���"�M�'?� ©��7K!�DN�l�v-g�������\5!�$�-o��jt(U�d���2��k!���V����IZ^��ځK�1!��]&ͱvÛ�y0�-H�*��t!�$�q��$�afϬ7ׂ��Љ�e!�}���`%ËuQ�0�E(� FN!򤐮���i��k��2�i8�!��=x�	�3�K^F,E�Gk!�$R@���T#�Z�����爐��	4��UQ��Q�)�'��|Y�b�a��5�Qi�j%Jчȓo'��w��k��$�󫄗/oBm�f�>Avg�-ZԐ�N~�=��E��T���k��6{BŀtAAm؟,��K�"ͤɢ������6ǐ�U�A���Z-yTx���	�H!Ӷ�
.�:�:OEy}N#?�ʙ�\d��T	՘����Y�(+G�ԥE��x�g�=H4.C�ɺD����R�)Kb�@�i
)j�6�Kcv`9ңIYFE���O3�1 �I�la�4�Q�'?0 @�'��4Ri�\�]�QF���K�SyR�̹'Hzta�+���.C��<9f'Eq� �1�+1`=a"GY�X%K*�7^��t�$L-qxU��EV�2��d�5�'��@��i }��Y�B�J�Ix8c��D��M��;���S��O�Bm�soT�M�Ԡ���O	I����
�'|���R��ر���f��O�t�v N�����W>��"��!�T�sc]��B It�"D������;h(�!rdTr�Uq�+C�����	���WG�3�	:oPQ�Vc�-+�@����аj�B�I:n
T� �����I�*C���G��8aqϽ.�����K~p5���3<O>�ꒉK4r����ը�x'�M+��'&�]�C�-,��=`��1c:����S:��Z�m�CH<1rd��f3f��05+�px�j�'dT	�,�24��`��i��UD��Rq/l\�H�����O쓁,���T�~�t�[�&��+��a�^禕�Py_*�Q[.��S��M��*I�[�z% g��}�(��_"������B���(��Iu���pg�i���Eb���3�O���e��<C!�8S�<O���I^��\3P/�	E� �@��b���C AL�� �>AD��k��@vI��m �듌�9>�@)���ݙOl���	�/��HS�סro2�9��^�I�3g���u)�G2yEz��\Q��E�ƒ����a�,'��9��NB!�Q����ט'#�R`��Q�Z"�k|#���Ӽ)�r�˟q�\7-��l,B��#�5FW*�S��M+�n�u;��f!�1c9��2�����^�;�ȁ����>�)�0Q��cy�-�E���r�˺>9�a؟y�h��	3�(O�9��
:Np܁w��ݖ�����+�.`sJ��{-B�!툞o��#?)T��R?��K���8=�� ��]���&�&_~�<	�e��?��#�l���-�<���'d3>D8�-J [
�8�B�PL%G|�,F�	��Mp���*�"���	_�6��0�ĭɛVE�3^6�� �������ٖQAF�\c����QkT�k�u���	mL��2�'�~(�T�ԧ*����iЃ_ *��`OǃM�F}��O[*��e R����ST�'J��Y�J�g�� gN�H�� C��̞$��y�O�T�u�#m�!Q傖nW8��E������+��P*`�V�^�����܂[� 	��Pdib��$�^��a���p� .�.x�բ7��r�'>�*�󨞧v��@�7�;*��p��:���iSۊ3q���M7'�R�lZ�1j>P3��Q~����${����2t��c�-}��ТT����vJP4иpAs�ˇ��>Q3'˅�z%���T���11��9c���#��9�.�	5��c�*�<6 ����
R�� b
��J�f5����+�6�=��b7<���1�r� s3'
-N,FEc����Q��.Tl�5˽�D��(��K��.0�.��A��^��p��86���z��C*f����ȱ)�¸O�~����N�cò�C�̄�t`��"O�I`Ђ�;K<�*gJֳ:�
)�0OJ���$��v�~���Q}��$�@�S�|�Z,ae�����g�v�T�>��>���<uz��"��I>��%�@��[[���cn�w˘B�ɵt�F�s&�XviA�&�Dad�=�Q��4R�ҝ!$	6�ӏi��0��̦�B5�EKO,I]FB�>xBak�Q�p��B��J5}�I�'�!wa�h?� ������ѝq����4���;f�8c�A5:�"����J���B䉗C��T3�ɞ�-��u���nx1���1���"L8�?a�n�A��\;�'-��U�?��7~������[�a�J "{-!�����'P���@�bR�38��Z�f�h�+/,�@��y��)M�R���x�{r��L��e��%S���	� ��0>�5�N� �HD��$4~�y�ChD3:���5L۶q:��c��;�Jt`#�\ǰ��dʇo���PO֭S�R)��c����D���ܗ	�n%!��^��z"��;!�Q�Э�?����&J���:��'�Ûx\`C�I*Q�|���m��t��]0g�ͫ1z�:U��<i�b�g��v�д2�P�V�h����9��}��vne�'*Y-@�1I�"Oցx1��e��5��J�@[�H6)]	Y�i6I����ht% g�󩙅f���{B�\r[����;8.,◣�8�0>�1��ұ�V��Ua�m�(k��t�ǫ�2j�`�8%�\ܚ��VON%~������=eO��I&�RA�ְ	2�G�AV��e�6x͒��㬜�/�2�qC��Y��d���	"2u:!S��L!q)Q� Q�)��B�& kr���痯]4ư2c��9|Ba"���M{v���L*14�ܘ�ԧnz����:� pX�B�p��p��̥���q"O�xfC��=
&P�6���n�t�4*
�a6����nQڠ��`ȧO��.�+��4��B ͽE
%	7��t5�9��'��=��n�8͂��d��O6�򱡛�4x��F��}�
 ��'�9c�g0m�a|��2$�Z�q�k˕w�(V�ل��'(�	(��_�̚tk�ɮ,U^�	�B��d���,5j%beK[=%P�"U��0B�I�n�FhQf��!Wy��QPR`�ب�担`�z��^�@(�A�k̹j�N`�}��6����ǫ1 �X��n�"��Ҡ"O����!��X�3��jb�Q�"�	Muz H��	'?�~$�FF�$/D�bp�)�I�_<ܡӁ%]�n�J`CK�\���M6Cx@9�C�
|�t�� �Ш���+J�$�7��6E�a&��/��a�R�ː}&���.A�%qN�>^)"�F_�O
�
db�O�R���D;;�D@Q+D*i��'�%�C� 6:�ID�pd���&�l$��kIDX���p͋�K��dpBiJ���e�ؤ ��ˍ#�`4����1���u!_l�����6;$���"OLP�3��a���A�T/a�mC�+��?�2P#�	�xP�*VA�5b��Ƀ�`���(d�Z�^�r�G6l�|1�p�n0rc�X�]l�?�K�n��)�A��Z,"���CzU� *+6Xbl*&��<z��&�M�'3�8P�R�4\fhΓIE�d1E�ߜ$n`0
��_�p�Ez�H�'V��򠯎�47c�o�9��I6ئ@x�nQ
Ъ�=x�1OlY"�JN�{�j�H3 1ڧ��d�u����"������kV�hoZ�.���╠�p~ �U�j�"~nڶ�J�:�./�6`�@��?c<Ek酯'���'D�����Bb��<���Y	 � )pda?��MKh�'�ȁ"�
�?1eL�
Q�AAK	!��r�,R�J���ER�����#l�j�:v*D�.��S�K�9D2F!QER&��d��!�%�`��*�v�dǏbo����!G+��m�vf:����q��_�Q>��rf�2_P4�� 	�q�80��2�8sx�PT/�9,` G��BR�{K211��k�Ʃ9���"�y����m��t!0͔�
�'��vQN!�F)� ��	0�#|�O"q��O)V�
 ��#hl
���' ��5O3EƠ2'�ơu�6�)�΁[�z-�!�L+rC�{"۹XY��▊o��p�M�p=��b��j;�i�#'n���U�ݧh�8R�)Y>��n#D�(s��TlzN8� eE�xU�7�,��2_��*��Eb�O�2����٢9|%�q/R'H����	�'��MɄ�ş1Ŧ����\�|F�J	�'�e��
J��%Ò+O� @��'8>�X��c}v]��*��qS�'d�]�.��$PFDI�Q�ҽ��'������5U�d� ��H�?u Т�'FȔ#��?*�F�D��$\V�Q�'kHU�cEҝ.@��C�g(+G<A�'K�\C�Y#7" x��lϯ%oV@�'��b�Y!/��K��N?�����'Q�`a�LR�1#��j�v��'�4�s�Fށa�@e�傎1x�PA�'��Yq�h��Zآ�ͅ�xBj�!�'��lc���XI���bƤ$}��'x��D�J�l�;�aɕ(Y
���'��Z�e�V&G?+Rb��b-Ҭ�yb�=�dBB�#���q����y҈?yԈ�R�R�{���cB��y2�O�V��)	���:4�IC��=�y���iH:<$$�%,�d
�B��y��<d�����Eu��s���y�cL/1aD�X�À>_�2vN��y/�'&��,p�Û-E�4��ӷ�yrEO��N�P ����d��y㕵G�*t����3�` UA�`�<��]�[A������D�<i�$�-U:�U��@@�mB&Q[��
G�<���R#�]�R*ոT���4À_�<)��Y%�z�x�nF6T��pc�X�<��M(�&��2`#:<�r��U�<�a�,%6�1R��.Q��h��#�P�<)V�J]����+!r�8f'H�<�w��6��(��ί
���s�FO�<сD݉w�B��#�cd2C@n�<i�c��1φecW�ӱb������}�<iN�5�:PrR��eˈY�"�G�<1"h�k2>lI1��?4��#g}�<�N�_���cm�'�V�0��[t�<�e�/L=�v�9���0��x�<����oB&pb�N�_@���R�<� B��V�/؄�b�k�9�\i�"O���Q��7�����	n4�q"OL�D�U�r,z5�,Y8��"OBT�+�	�R(AFCy'6�ك"O���T�(����E�D.w��Ҵ"O�p+F�J����qnňx>��r"O6`�� @�jpX4^���6"O��9�?s��ʓ$F�v\����"O�(��E�=���Ѳ��#,gF1Q�"Ojq�ű3B�� fBd�"O�ͺ��ط5��DgC��'kr�A�"O�\ p��({�����\V Q��"OVuI֢M	C|������?p!L��"O�e���4| ��fS�QH��Q"O8e�G7i�F� ���tQ�5@�"O��yeN��Ubǭ<*XZ԰C"O�C���.0V̙�DJ.�ˠ"OH� 4b�����J�7IL����"O88�V�W���j0�w.d� "O�e��/��7�~pH�jϙm��4� "O>U0e�ߚ,~�Y'���tE�s"Oha��vzص��k�"��P�"O��%@�7-Yڥ§+�;J�@�1"O6�q�S2V���Diӭ
t�$x�"O^��0恗W<��!�g�Ր�"O~9+��D(�� bsa�+@а�P"O��I�3/� ��ג��53S"OT3r�}_d��UN������G"O�"t��<����$�;�4�3"O�
�3GD(�l������A�ߜ ����E�
�'.�=	hI��&?Y��%9H���i�
�\%���%8X����Xa�d�>��c��"c$���L�4n��	��9�)�?���P�N�p�L.]z�m	V	�@���?��\��y�O�(�(GL�;��
�ȃ2�&�8��$>�S�$	�,����+A�S�`I���3��'R�I|>�5���'ϲ�BQ	t6�qU&??��O
b��'��ת8H�`%�E�e4l���F�r���<ٰ-�>E�4M*�����$vB�[W�����$F���	�_G`I��B;l�T��c�6i^�����d��yB�}�R��c�M��p��E˰m�B�Ie��ݠa/ӟr�$�3Ш[�%j�C�	�X�D9�N��6[���a^�k`C�	sj�d�@��
 `�2��Z�`
�C�	������8��\I!���w�C�� ��1�C6��D T�@
c���INܓ�0|�F
i����'5f\R&l�<Q�I<�yb�ijD��Z6L�?�Cs��;k��� ���nb��Qu�c���`Gm�48�m�0��4����0��ħ{@�<��ǆ!{.�K�˽�虰���}}n�Ē?t��؃ш�I>��JD�@�p�,]���V��$�vLp5 V9n��@/l�H���O��A˱K8|�Ř "K�m:4��_4�V���Xxis��Ih�Lܧ|�Ji5�$j�Z��4]-ЀÇ>O,M���� �E��"Mx>]�d�P�5�P�д�\�o�D��Ê~ӎ���U���dě�y����4{�񖭓6���!AϿV�.I��@>�����=�)�$j��P�-҃���`��GdK���`��@Zay���M߬9ۅdӚW�ꈘ����y2���pܣq�A@}Vl*6�ɚ�y�@�)cb��Y�JM�>���b�d�)�y�ƞNhr�.Ӓ;L��!�ʽ�y"�D�<��"� ��=8D�\�yRK�' ax�LT	Ꜩ����y��<	H���A��RB�5g�Y$�Pyb"�..�`�̆�z��P%�g�<�Tl��q9rHS�mTz�MХ"M�<��G��h����
?�VX��Ec�<� :1��	M�J>p��Aƅ��0�"O��hV,'(�����*O��R�"O
���͈:����to��{0���"Op�:�¯~��z�g�	;�	�"O���ѹ$HИ ���p�&ճ�"O�L��/�	IU�܁rIFF��j�"O��qB�c��-��GA�I�f���"O�1;6�<(�$٪����N�� "O��i�OC<����d�� �h|9w"O�1q��"����ܻ�"���"Ob�W�̙R��D��T68g$�"�"O6�Y#��q����a�N,>�FI�3"O�U�p�F�9��1�Lߊ? b&"O�ӊՏB����R �P��"O�`��_l����	ފ��� T"O"��&��$��؂5�;3�4I�r"Oʍ���A�
=j��p3�M�d"O6�cv�L��Yq5�*b���p"O�[��	z��e�Ţ�0iW"OqA�~,���J�!����"O���SK�E�$��J
�*�6t�b"O,�*�D(S�T�)B*�e���Y7"O���b�Шy�)y7I�Bk^�ٵ"O��0� C�<�S���F�ԉ�"Op�B�Bq�,[���f̄��%"OPm�E���:r'B#i��USV�:�y�KL�J`a�̡gHr�rb B#�y��N \�`43�DH�^o"��4��y�bP.�(�g	C:(��bB#�y��q &QC�XE�x8d���y�"F<u,u(#��.����:�yB�R&e� }��O�"��q��+���y�hR�u��hrb�2��P-T�q��'`��Bd�-5��@���ˠ�	�'�XЁ�ȉ	:��1��͘�a��'&tؘT���8�}�A(M�A
�'Xu�4�$X<TJ��?;`|�	�'�X@���T}�y3�'��*�M�	�'LP9ЅG�Mi��B2Ϟ.TR�Qh�'�^�)��!~�d0���TX^=9�'�e�FO�����U0y~M�
�'䐤��Nb�2���Ɗ�4��'����4���A��S�q��1��'V�*A� +ypj�g�H�8�'>�%�Q�]�~3J(�������H�'� 1V��51l"�z K�\�q�'"������t��áB	���C�'^�%�G�գT���BaߋU�t���'�t����4_!�a�`@ƚ>rd�`�'�p�3�)6�I�O�b���"�"O���4�C%2�L ����3wfh�"O��b�*�*GԄP��(Ҕ_���"O������8)ˢY�@�ג]Y�J#"OX0 w�^j�Œ��ֹw�~a"Q"O^A��Ů�H�X�����uBw"OtM�&N����l
%#��W��c5"O$}�p�N�ԩ
�^=k��� "O��ȃJW%;S��E H�`Ҡ,*f"O�E�%��8`E��YE��$@f&H�#"O�MBReN>H�%��);R� �"O��c��Z97�1���˾r">L�"O����-Ģ&Z� �s�*4	��ZG"Ov�٧�[�t�@���L�^���h�"O.�����|�ޘjWG��>��1"O� �h�HH��.}0�'@�.�^���"OTi�_�'����� N�M{fU��"O�����Q6��`/3��ae"O�({��Z  ��/I�˘��"OR�%D;<;��al�\����"O������d��c����5����&"O�͸�iԃ4�-zv���x����"Op͹�,�E~��3L�;A��%��"O,m��B�*g8�`��"Ҽ�"O��r�'��D.�L&%P-$�t�D"O�5 �ݛew��n�9,> ��"O�ŀ�σm6�̭"\�j�H�M�V�<1�� as�5�".h|m�v��Q�<)�ON��`�Ye�*P��B1KP�<�/�>cT���	��s�@�G�<i�,P�l�
��V�F�Y���K�)	L�<)$���EWp�ؐkC�K𠔳2GS\�<W�¢q���1���<)���j�V�<Q��.V� P�RF�.d�nLb�&IP�<��.9�ؐ�/G������e�<!�$�4V��U��%؞O[$�B��\y�<	t@�,��!35�I�`Ȓ7�j�<�S�O�Z�&�� Q숕ʡęi�<��wҌ��#�@�gP����n�<ɥh�<0!�I4��5�n�P`�g�<!�e����ɶ�\��-"�ǔb�<���T�yt>Hs�lA0�9��^�<���6%��$KRD_���BZ�<i�$ D܈Fb�5	�AYp�F_�<9P�9�X%��t"*Uy�o�P�<9D��F ���ǈ^(����P�<��Nɬ ~��$	_�W�V�($�I�<qA�L�^�XA�e�J"�l�ȣ��D�<Y�O=rb�[㮎r��`�CJ�<1����&�
�ʆX^��I`�@F�<��-�02�Z�rT[�PP	� �<��D�
1���a��g�@��&T_�<Y5�Ѓ�,ڕNа4�z�8�*�A�<V�Z'���R�圡,�LQ��� t�<��m�b�n��#��J��)A�z�<yC�+I��b���1��O�<11%�-`s�@��E_2���@�I�<9F��-4�X�2��qpN0���_�<��+^ج(�+p�VIj@Y�<�p�34�R�f��2��iBS�<�0)'p<��j���h� #�V�<A��a��ׄ�5E�<��7(�F�<1v��[�Xy �#��R(*G�F�<Yc²��E���O�-�*�aC�F�<�CDT
M��D g�ц:Q�T���K�<!r�U,��j�f+�r�	w(l�<y��%D�@��"ţg
z)�B��h�<�paQ�F��I����.3�Lh��b�<���U9&�~��wo�#N4�j�C�<�Q�k0YA�ED%J*F-�j�C�<����{d�}hQ�� E5�T1��A�<)P��h��sd�6t��"H�<	T@U�!c�m�An�:wN�A!��N�<q@�t#R	���U/Og ���M�<	�#��s�&���qu:L���H�<I�LJ'^'���"B-*��2��A�<�B��+��\AR`C]���r��<�`��:`ᩆ��Y�f��*�}�<��EȲm�~� �S�6�j�mKz�<� z��vۮ&[���U�>A��Iiw"O��{�E� ��A֊�m��y�'"O���`���ji� �Ui�2S��)@"O"ݡRIۤS�+���9g+��j�"O^���Gҧ$�2�)�a�%r��"O�i�/� ��AA�����$"Oةq"�"X�2����7f���"O�]���2s
pe�f�/�\j�"On<YèJ�y#�%�� �� ���"O��*�e��P���eƏ�D�Q�s"O�Q��
��@���dĩW�4��"O��P 
�3*�d£#�^��L�5"O6X9���f��{���8S�1C�"ON����� �\�bT* ,Dpx�"O��0q*O��D�js6<qd"O0�����*��h0&Bl�L��d"O�Px`�R�Y��:p�L)h�p3"O��	'R�2j|��Ae܆*���"O��#�̓>jLiPs�ϕ *p�p�"O�(��΅I����B��;��Xu"ODIH4g�(4�@���(*�$��"O-�R
��~h����c�h��%"O�-q�(N�*�,p���T7�]��"O^H+���$��9���\.-Sh��3"O� �!d4��(s��kX�U��"O��!����\�ҍ�PV8B�1�b"OnЈ2晨Rʦ9A�@�;R��"O�,��+�:4�dL[`M��yq"Oby�de̤D|(���/�����"�"OJ��m��n|�0!��=z��q��"O���g�"���IfR�"Ox�B�,�+y�xd��3Sj��v"O�̂�K�t�	�������q"O���Kİy�T�����l)v"O����	TP�CR;1�xH� "O�l��G��YL��DB�z���+U"O�8k+FE~͓2/�~*��c"O�4��@q%� ��< �4Y!c"O��{A��W$�@A��07���"O0X��Ĥx��h�S/��Ҭ�"OF��`N-r�|2"�
����"O��Q�F�<0�h|�%&�.w��@�2"O���X�^��c���6R�ҹJ�"Oh�! 
"j���I,Or��&"O�a!uƕ�o�N�q2G�g_B4R�"OX���%�uQC��T�O�)s�"O\����>d��e)~@��6"O|]���4]ĉ�J)Z�F�Q"O�DHB#R&y�����(!!Ȭ��u"O� 2�R�I���s�|ءt"O\�s0ぴ��M��--"�4,@"OܙI$�
rp��[�fޛC�(8{�"O����U�,Ǭ0�6F����1K�"O��(2�d��iwb�0�J��7"O��j���Y.����@�m<���"O|lY�@�;S�)��	�Pc��ѣ"O�=����E�[�nϥ�@b*O�`��Ŕ)K*�=����.s�B���'�<<�q�94$�91�M�p�PT���۞<f*�oZ��n���M�'r�.� ��?A��MsY�<���A4�d�«G��,%a󈝏|{	��3Ҹd
S(�?Y�OW��@��<��"Iw�h��#�r�l�Е��IXq�'��mW|���g`���;�u�g%�iEļ7�ْ3>���fX,1��Y;p�"�'L�6-�O�=c��Y�(�+�e�^��P��%3v����^�?َR���&�ıj7� X�"�j��ڈ.5"�H�۴*2�����x6� \�2h��h��Q�2�\̲�����,�IR	"\N�I�h���D�ZwT�'���O�u���H1� K綔R�U�<m ���
 &�����1�iȓ!�"ψO��Qƒ�LƠ�AٟO�R	 �YKg��ڴ�S�x]�O[��Mc�/��a�D��}��+�p��E�4�y�Vo���Ms%c^ڟ,�I��ē�?����ēzrj����F�PlZL�0A®F�X��?i��?��H�`���)OX�d�HR��d��kf�0�O��l��?i�'d)q�/d�27M�[���@U�]����)T&�Zt��؟��	!L�Ĵ��ԟ�	�"G &{B�#��5yR@`��"|���%�L�K#"�+g�ȭ®�����W�)�܊�G #(��d�H�'0��(��G�&��0�<w�D��Q���N���
��	�\���O��fL+{�n�����U�ص�
@���I����	F�	�'>�
`K;	�I�7�N%�@��
7D� ��o�?S)��i!b mx��;�F�Z��
e�"�DTߦ�Y��,�Mk��?��
2��$	��D�`�83��١pF0aZHA���?9��&����޹6�`D��"4��	h���?	�;[Ѥ�X�F�b��� �a1 j��>Q�� m�,����_�~:���0��<M�1�[(iJ�P���P���*8:�8�$\��+9:��ɢ�M�ֲi����䣟^���bP�Hpv%
iz����$�O�V�hMy��$\��@�w��Cs�$��	��M���ip�	�Q�q05Ð�䝛� �[�z�^�[[���'q���D��9 ��'O2�i������c�j-��E�n�H�Eʂ�M<�9�	��\4׍̈́x��)�|��'=���	�c%���{�R�"I__�
�:�D�f����̉>�(����YKʨ8���I}މ��$-�)���M�n�]��ǜ�?��-V��'5��G��O����@Z�h4|��8S��T2��K�x��e}"o�F�D��ȋ�eS��B�I��'7�\㦡'�Лeߟ�6�ӷS�N؂w.��Z���F�U0N�<���~�.�RQ���4���\�������O�7m��d��6�S�d!���4M��I[>�١hJ�Z�aJV��|�恡�eM*��ْ�/
���KV69Sv�@ud��B`h��o5�`�3�
�f$�֝����[7�U�.̥O���%"S��
� M� pHnP0e��\#2���!�M�$�i�_���ش��^'I�2�O�4��i���|L왆ȓ{�>e rI���)� <kN1�wJp�(�O�}b�O��'��I&H�� �  ��   f  N  �     �+  ]7  �B  FL  1V  %b  Bj  �p  �v  *}  k�  ��  �  7�  ~�  ��  �  E�  ��  ˻  �  P�  ��  ��  X�  q�  H�  ��  ��  6   ` � �" �(  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3�����M[��хJ��x��#��+�$a��)i�<)T.�o��QՌ\�@��wga�<���4x�����KyK��jBD�^�<1�T���㕧]�_�D�R�(���D{��)R4i��	�`��>wܰ=D��#/$�B�	?~Dr<��E�T���W�T4@��4y�\Fz��HR�K�  *��[�_H(�"�J)�y�X���!�WDٚh�"K��y����<��mC�"f�d��C3�HOУ=�O�z�y�-ˁy��ey������ �'�ڄ����H�J���+� �.@)�4��>R��uG�s�~�{v"@�O:��ǭKS��H "O��*b�<��25cݾt�T�9��R��?�{����鳦
"�|�	u$C�_�D�s�/D�h!&Jo@����ꋻJu��o�n@a���s� �1E�Yp�r}�Ąʇ+=rI%"Oz�3`��U?���P4!�p��OL��DM�y�MX� �9�H%
08W�}R���@G�KbF �2�W�'�&Ö.D�Dò��RX����F@��\t��!8��hO�%g���X��}�a�Æl�nC�ɸ9�K&����Q;!&ՒyDc�اO�ME�ĥ�D)�d��.�"_k�ْ�mV��y�(��ȹ�E�V��%�DzrH-�MS��O�A�r�lڧ��I)��w�$,��"�	D\фɟ-<Q��c�'+d��v��gG�0���8-�� �(Л�8O>O�A�Ϙ'H`so.%�(��2�J5/r��O��&���}�Tm�Ot!�@HA2%N�k�%�>c����"��(x2C�	�f�.HH�kB�.�2E#B�3B,B�I�q�����	\L^�s����C�I%�e�g���Q� Q���yb#=�}r���q.Y3Pj-��΁�y
� �����;BL�Jp��|��L�c"ORm2iQ-���	֮�9�~E���TEy��d�OH��fiP3)O\�C�GܲY�80 ��i����)lUL�Ŏ�Tf�)A(��dc�Α���~�A���Վ!��`G��|�Ħ�S(<۴Fx~���
�
�8� ���D[��|��$\O�;s�	�&�J�Z�OМB)z@���'бO�ݒ�C": �|h#�	�I*U[�"O��b�A\�H6�mk�!�9I�H bR�x��)�� sb�]���B��k��?�b6,������ 	Oj-А
ܑ_��xar(&D�؊���#~���[��E^��6�$D�D���"�Ԉ��-=*�p�Yf(#D����˛,d怜�Wgֲ?B���3� D����AL1~p�h��4����/+D�����f��,~ucF-٪&
tB䉤=kʀ��_�ؤ��R�B�I*[!.@�.�#I��K�e�+٠B䉪!�nH01�̟]w����GL#O�n��D(7�D�T}��$�41�ȓ	�]�f�%h0�)���d3H���q�����fɯ�T��1����\��a�z�	d�M%:�H��%P=+��=��4>ay�들��L�'N�@Zh	��ƀ�yrD�VÆu��ت0�r̰W�ͷ�p<!��䍰�����Ar�KY�u^�	��M�O��a6[���h��@AՌ�����ȓm7FI�5 �?���c��Z���I�9��I[�j�1�c�#X_`�P�D�>�C䉟z�,,��ˀ�G4��U�)!{z�O<0��'��ı<qI>!�N�_ÈQ����S^�����t���'�6�KG�TT*D3/��ц	xY��؟�'��>�� Q�\��q�D�l��9F��#<ش����O�hiE��(b��[t!�� �
�O�Q�R��v�	���#����g�>��4��$4��L~���5��tu���`�9�N�'�yraݛ_�$a��Õ�UqB���I�����?i7e+�
��ĩ>�6�B+;j�+�M��=�P�h��Q�<Y�[7v�RA�U�&qð� S��Ny"�'�������;%�p[T��	j����'%x!�GJ@*Xmh��[
�����'�b��Ƌ��
fFMQ�I�SVV��O<�����F!+�l1��a�:�t�U*��P�b����
ۓ%���Ԫ�?��
�IB�L�xO<��D��P��� b��؂v�}+�)rf��O�C�I�1�rUPEԕ<����'��'�B䉥=>��тQ:�r����KN�lB�I���S�#R/.j��è_5j
�C��&	�^�B&Y7�D0 �#� ]�C�ɃJ`�gJ��)J�k�:6&�C�	"6�0lOA9y_��ئ-B��xC�ɫ&�j,{5IX�:F>|�%M�0�C�	�a��M��|�� @	͓O"��hOQ>��	!o�f<yF�7Q�� �Z����8ړ	�������Wu�X�$�pȄȓ$fE�t隦hb�ʀ��0�T��ȓ
nR�APs�&�R1��"_% i�ȓ0��ƅP�,FΨ8�$T���'����'�2��+�Iʚ1y��=�VI��'R\Lfa�	#RL�U�_��t��"E9�S��?�r��4�X���^.]��LP��S�<�V#�7tVE��G�/1�C�v�<y�ʇ:%Y�H&��ƪ�oVq8��'�\4o@}6�0��U3-_�A� 8D�� ����$�f �ma��m@a�u"O���dW� `vBQ�D!Jԭw�<�A�	S%��Y��	i�ʥ��Ky؞0�=��kIE7����F"�~\h�'�v�<����na �`B��.��$ f��M}Bb-�O~Y��͍DWP(�T)
c��D[v�'��6�zlЉh�$�B�9Ъ�DyR�'Ԕ��cIH^v|��ҏ:y:<X���;�������� ��[F��~>M�ȓt$�IP�X�&�� ����ze���I9�?y�}��)�&;	�	aYNj�h���#*B�ɕ\4���t�S{��iRg횄wV O�����)C�kT���!�����lѶ ��*O�9�� yp�,�7&S-<91�'��C���=�Af��2-���0��D$�''�tx�TB��D�V��A�(��l�'h.�[\�ɻ�&��o�ƥ�ϓ�O�Q�A���S��a��g� � �d"O���I M�R�	�FͧS�&4z$"OrD�SK�LP��Ks�Q9,�F�P��'G���D�����$ԲKN��cb�#d�HC䉦�\] rfμ6����*4F�<�,O�#}2Vo��h������%=:ux��P�<��Eϣ#4J��DZ�UF(���<)����Q�:�j�ʗ'$�2m;��2_�C�ɚI�$�x' �d(Qc�]'g��C�I�c��,[EÕq��HA捛�`NB䉜
q5�ӋY���Ë���C䉣"Q��;�.�97�4��OI��b����'�a�Tn�:��mu-.C9����
��y�ܚSTlM��-��+��Ĺe� 	�O����p2�-;��O�Q+�5������!�DG+S�*\0�EP0_�p餀�9S!��ڼ�8U�T��*c���0f���!��ȉ8�r���l�"N�����$�!��jf.	��

�7?X������!�D�@�.� N�#b���.[�`!�D�X�z���� q0u�g�_ 7h!�'H7^L�
2'����,Oy9!���Q��m�>h�^�0�k)�!�D�<[��h�A	�Ẽ��k�?C�!��A6|D�%[�*�29�.Xá�� }�!��ػvvl��ē����,I�!���!u��(�b}S�AA.:;�C�IA���7Ec�I�" �h�C�Ɇ;���mW�h� `&-�$hC�d�:��Q��S�
l(�]�7`C�	;7�8ɑ��L)XK�(u�B䉟j��AG���Mt�5��ڮB�I����#���d�x�9��G#-j�B�	�	AF���j\��hH꧆�
�B�	�x�YYQA���{��KvR�B�Ɋ6��Mׇ�u�� ��"�2,B�ɝF����a�'њq�=�B�7,�&���/Q�%�����9(q�C�I�V~K�.Ń0x����OE+��C� ����k 
_�������)U.B�=	�b�H��)x�(���A�=�B�I+%��i����M�dt@�c�>j�C�I�%O&8��̗��>pR`'_�MYvC�I+66%Ӣ@�*6�x�($h���"C��1<=�@**/W$����w$B�	�__��Xw��:�����^�uB��89�`�pV��e朒���65��C�)� :�I�Ç:^X�hq@��6!�� �"O0�2�>Pp�@���^=���2"O�5��6#�}�2ĕ9]�i�%"O��SM�6��d+W㏴�9p�"OR`��N�iΡ��ʘ�S@�'�B�'S��'VB�'���'���'��T�4�ހ3�Ts�Ѳ\�,�*��'�2�'�'Sb�'��'���'�$Eg����x`� ¶�X��'y��'��'�"�'�"�'���'KdP���Inz� �`H�o>x����'���'��'���'=�'��'T�HR����D����2B�"����'���':��'"b�'��'��'{�9J�$L�^m8�[P�s�̐f�'MR�'���'F��'C�'���'6�ty�jKW�����돠l���G�'�b�'���'<r�'���'P��'���u�B&<4�$�F8qr����'Ib�'�R�'t��'2�'&�'��QE�F9T��SAʴ�ݩ@�'�B�'�B�'���'���'���''<u�.Մר��cAķvK`�Ba�'���'�2�'�B�'.��'���'�Ѡ����F�N׫%t!���'���'���'Jb�'���'r�'�\�9 �X%GϚq���ʷ6�Иe�'�"�'�r�'���'���'���'����L�|^��BLQ�	R��'>2�'��'���'��-l�8�D�O�-��Ϡn�5J��ٷU��M���ry��'��)�3?���'��)����<*�]�r$���J3}2�d�v��s����&dr��$�@�%:A��99rh�����ЃK��m�'��I��?���p�fƜ��$�8�oƗ<o�xp�D�O�ʓ�h�� K%�́�Xq���,5N��  ��}9��*���MϻV� "�	*Gf������	���j��?	�'�)�2�f!l�<!�'���&-���$�)�%C�<��']������hO��O����A�Rc��B�k*t��2Oʓ��.���&�J�y�4��Vb�'Bt��M�+r^u��r!�>���?!�'�ɦ`P���h�p ��H�MD�t����?�!��<���|�1��O����W�쑉T凔*0��I���J�r-O���?E��'�`��疍Gc�����Ԛe�f\C�'*67m���ɤ�M[��O�6�2�k�'k���!�ᜟWH�ș'���'@��+���� ̧G+���h�X�J��C���c��πu3��N>Q-O1�1Ol��V��
Ѩ���΀��TH@R����4"��{���?Q���O���C�1v���c�`�z��p�N�>9���?QO>�|bѤ�$$� �ҥJG�ci؃2��!��񦥓/O��7O��~��|�W�s �ˆb���E<u����ae5�OBoZ3R�I,�p�Wh�,`mP�K��[!i:�I4�Mۍ�>����?��5�usq ԏ �E��(�:��#R��MC�O�:��χ�R��/����:h��`��\�l�����D04�P?Od���؟ ����Ŋ30�ȐӫC�#��˓�?��i-rL�̟,�nZV�	3P��p�0*�B
�qZw�,��8'���	̟��v�8�nZi~Zw���,�J\�g{:d�v��4�2��G�Iuy��DŇ(�CW�ϭJ��U�u	A*GT�d)�4�`���?���	���
A@C�Qߢ�JS�[L�	���D�O���0��?��E���^�g�$U�#I�^�|M������*O���~�|B��/T��
ñr��D�Z�9B�'���'o�O����I��M{2!�3L*� �(NA��9j���2A�����?	�i�2X���I���d�OT!2�E�5�rh��˃3yt�r��O�$M�r�h7�e���	�jE���֟~�){6}��ңe TB�PYEfQ͓��$�O�$�O���O$�$�|���b� Kp��AG놌�`)L�nZ�I6��I៼�	�?A�����I�杧~/�Q�oR8$����1��G;^y�	U�Iܟ�S����ɖ '&(l�<��lG(������'�E�,Q�<����
Pp��R�W����2�KI4(�ba�C�ս �B�I�
])U����dc�-V�~��C�ۙ�j8QҀּD*ި�ElU:b-H�/�q�=��e�7j��r��ԇ:纘Q�ۦhrn����(�깈@Z	m���s� Ce"�Z������6*P>:��0X���*���  �X�a�:��I�SGd}����-k6�b-͍3��(A�c�
�r�z��A��
���jFx�����J�*�(� &e�9����3r���Y3N�h���a���F��a�'H��nqŬA�$PTI�g*�F���t��Ol���O8�B��Ň=�0�%+��V�x5�������	n�I����I�/gH��=��Ҳ3c�|铊�Xq�����1�I֟�'�
�*aY>�Iٟ��S�e�^0��E7D H�� �(��BJ<���?Iwm�������A&�V�3�4.�tyH ��?D�R�@��Bɟ��Iɟ��	�?��5vk�9X��.e�XA�N�Z�n]o�����I4g5��?�~rN�U��r0���@e mPq����䢟����	埈�	�?ŗ'�b�'Aډ;��ԈG X����u�|f/w�J��2,�OJ�O>�	&Rp�@k�D&�H���J� SHKܴ�?I���?qb�ڀ���O����O��I�{26�١J��w�2��R�I>��b� ��I+���@������ �d�ݪ���@�_���ԵiG�e^"{<�	�����p$�֘�=���Tk1N~*�����o5��%��������$�O�$�O,˓z��#EROL���a�
�8r,����O����O�O����O6pᤪ�?o� ����i�4�V
��t�1O��D�O��$�<y��ʫ���Ɋ�,�`!��Rh\�僱�M;���?������?��q���p�YN��)�/7�4�;f	�;_��`P�x�	����	Ey")է}��ğT��S�/c�A�#�>r��2͒
�M#��䓕?)������{BB����?�ԚTσ�ڼ7�O��ħ<��*�|���Ο����?� +�Wt�9�F)�4�N`kU�S��ē�?���E��`�bןvX�'�N"`����C(�D�7�i�剷;������I���IyZc�2���'�\�X��oS����8ݴ�?���kP������O�5J��8`�Y8����J�
}n�q*�@�I,�	�����Ly��'�r��P���S�Ĝ�?���ؒ��Lm&7�+w��"|���@�8�#B	�Q�E��BRt�9���i}r�'��M ���h�I֟����t��p��^܊��Gz�h�>�Ə���䓖?I���?��5��cJ(�rݚT�߾h���'�p�P�+:�4���D�O$˓5&�����P�� �Wi�/�l"�i �m�=q�rR��I��8��IyR�K�2c�U#5�$�$�:Kp���1
:��Ob�$�O���?��OZB�:������z��W��ڴ�?�H>y��?�(O�L�Vo��|zW���F) �P�N�%)���FTH}2�'#�'������O��B֛,.LdJPaB�d��kq��4O2��O�P�r+q�������	��kB��G�q�f`��4�?A����$�O���6.���|z�+�INl����9��8�W�C�a����'V�P��yQ���ħ�?	��3�ݔ5@4�`bW�x���k�ަ��'���'"i�7�'��Oq�\cxj��F��C�9�S�4�(�ش��W�`���l�����O��I�L~"��(Y����djؙ:ꔡ�qL�M��?!Q.Z��?	S?��I�?���M�ʀ)X����L
�_d�0@�Ǧ��AC��M����?	����%�x��56� 1Rp�@��!�l�I��۔�M˕F��?9��?����.��$�O.x�ċ�J8�L�E��c��z�������џ(���K��N<ͧ�?i���E�_wP��X�J*"�@
Sd���M����?A��b!���4\?��O���O��� ��Xg����(߭ Ɛ4�iCR�G}p剦���0��~A��kR�SP�E0��)]T
1��O4�P�]jj1O��Ļ<i�2@�ZRH�&MF[u�X;S��h���"��$�O\�d,��럈�I09���P�E������%윒�쒮U�b����byb�'+ \�cڟ�ܨ���!������>s38��U�i�b�'5�O����O �q���Dț�v�M�!���@�D�*����x"�'l����ƥDj��'�0ً�h�;�!����_I�;�pӘ�l�I��F	i��OD�����{I1V�Ӻ4
�pIŶi�bQ���I'�Rx�O���'��\c���"o�f���`�ɍp�|��K<����?駋��n���<�O��ydO�m�\T��M޺d{�y�O*�$-�|�D�O���O*��<��T��8',�C��$��osJMm�ޟ��'��`���DBД�\QI�iU<Fi��Ч��M;���?y��?1����(O����J�IH��j"� �"Ȟt��9�O�����)�ܟ�I�ȸ1zԲ�K]^�؅�̥�M��?���*͊����x�O��'��b&ǥ=��Acf�_^�qdi{Ӛ���O���^�Y�pm��yB�'���'ar|J�Z�&;KƆ^�H�8v(�G��V�'�ʵ�P3�4����O��(ֆ����>6��I�L��$�i�"��4]�R�|��'�B[� xq D �^���>� ���d+�T��I<y���?Y������O��$�I�V P��ܓ7h��H!5��(���O��Ot���O�˓zܱbG2�.S���Ls��=	p(���P�����@�	^y2�'��a֦FU��N;e!�xv%�.�JL�oK�qT6��?���?�*O�=�ჀI�S	?6~�jF�"O�.t� ��� �М��4�?A�����O��$�0^f�d8��B�[��	"`	�h�ځ !�Ms��?i���?	�朇b��6�'E��'���㖧4�� ����CIb�p�K�=�6�O���?����|:���4���gZ�Y�rD0Püy�Č
���#�M(O,C�&�ЦI�	@���?��O�;}=�`!��c��@��O�؛��'!"HQ��yґ|R��6
U��(搓 �*���Z)V��o��6��Od���O���X}�[���RYt�,A�l�Z�Y��ʊ2�M����<�����)����0@����$�q�-�C~��arȎ=�M���?	�nz�q�U���'���O��	u��/-��0sΝ�HTFU���dV�1O���O��Խ*�����A�����ߠA5~H#�iJ�#�z������O�ʓ�?�����(�B�9�l��c'ǈ	��7��Γ�?���?����?���?)D�}\��*HX�sL�XdF0� )�id�'���'��'���O(�D�7-ݼ5���އrƌ�Z�!S9C;��O����O�bӬ���|Ҁ�	�8�6�;� �y��D�87�&�㯍�M�B�P��i�r�'��'k2S�P�I)h���&��Q%��!�H�����!XV8К�4�?����?����?Y�w7θrƽi���'`D$J�T�p�Lꁈ�J0�x��e����O���<Y�2;J1�'�?��'��X;��.)��[�Z	:ƀ��ݴ�?q���?!��/����A�i�2�',2�O����U�UOp��ꅀ͝LȒ�ic�(��<I�d��Χ��$�|�	�L�uԘ.W�1�\& ���'��+L�$Vz6M�O ��O�������L�c�Be�&j>��Y$�C
d�h�'B(%k��'��i>q���kǎ�V�1� ;Zp�8B�i�	k�j����O�����X�'��I5v��][ ��?��S���T$�y�4_=��Γ�?.O��?%�	��@��0@�(5��4ץJ:*��x�4�?Y��?�"&�5j���hyB�'��$�%M��ⲡI�16���*^�/q���']�)q;��)����?���M���Q�502-a��Iz=j�c�i8��Ň �����Oʓ�?�1v�p���,o��<I ��%��!�']���'m�ڟ���ٟ��'�����M[8TQ@I����D�=z������O�˓�?���?	�/�7u�Ɇ�E8y@�#��ʘ��?����?�����9O�-x`+Z�|��a�0.����+�T��FI��'Q���ş\�I}\扱a���(�gɖJ,������́j�4�?��?������(UF�x�O�Zc���1�_�rP!�z�h.���]yR�'�2�'2^�C�'���O�ͻ�˧t�JM�Aà�z���i[��'7��tY�}��~��O���O8���5���	�C�B��',�')�"ɑ��I�<�O;�!t��3'��3���"�0qH�4��d�j�m�ʟ8�����S�����9��JO�(��eC�9J�K�i��'�*d��'���<�������>`�$DY<	ؠ�K�M���EM֛v�'
�'�$��>(O���g�@�[����茍'}�ԁ7�����" g���I^yR���O�$H�/�f�V�FCP�w�%�5� 榑���(�I�_:r��ܴ�?����?����?��6hd@�$@�y�u�f�H�k}�4�O��z71O��`�Ik2c�\q���a��9DV��W.@��5�ɰ66�	�O��?�+O����;�L\8P<x,3��_�q������i��`V��y�^���	ӟ���zy��=~)2�*�њS�0�
@NԪfo���M�>).O�D�<!���?y�u;�h@�[�+%�t�4AN8y��]�<����?����?����?��s�8Y6�iHĩL� 0 �(�gB�	Y� ��Ja�j���i��'��\�h�'/�t�s�0�s�bʤ^Kjx)E-�	,�B`3B�i,r�'���'G��'Y~̢��zӲ���OL�8�A��:�U�yd@�piM�'����'�2�'����Éd>���ӟ��
V��VT�t��T��@:�B���Mc���?����?��ą�T��F�'���'���\&p$��,۞~O�T�"�P� 6��Onʓ�?� �M�|����?�/��	��.��u��kU5E
���K"�M[��?��a� !���'B�'����O�R�� (^xӱ��0T�.d	w�@���?)p ]'�?����4���O�ؙ!@�Q�;=�-�B0dTꐑ�4\p�E�i��'o��OE�D�'?R�']R�JX�$��p� L�Wv:���e��T��?�i>c�$��.a{���H
����U�	j&	��4�?!��?�$.P&}����'�r�'����uG��j<����Uv��*��K=�M�K>�����<�O-b�'�"�Z1����S%9oVA��e!av���$�0.�&���	�&��X�1pm��,7��c��²_t��M/�������O\��2��Q<S�1��!$)) .>Ca��E�Q��?�-O��O��$�&vXЂ�݇d~,��E:3RΈQQ3O�˓�?���?I/Ox���Q�|��ՀWX��lW�0���pW�QT}��'��|��'���[��y�j �|d\U�F]�:�:��f&�+݊ꓠ?y��?�.Op����G�W��:�n'U>��$�8	� ���4�?aL>Y���?)�@��<)O��	g�PZ��PpBCS�ܳqmi���D�OL����sR����'��d�FD|�E'ڲn�r�C%.�� �\OF�d�O��c��O�O��8X�ke��<T�+Q���,6m�<i��<��̢~*���Ğ���Ѻ<�R��]�
��u� �bӸ�$�Ov�B �OƒO��xiBǢ(�hQ@UcԻU�Ѳi�e0��u��D�OJ����&���	;pƨ�s��o;z�#.-�(�:ٴ�H(̓��S�O��g�8��y3�ȅW&vE�@ꐱv�F6M�O����Opr�H쓬?y�'��ᤇ�<QR���7���}�&G���'JR�'��S\�6T�#"Њr~*�"É��*��7�O|y�ΐe��?�L>�1M\bܫ�휜P�2њ�a���T�'��a{�yr�'�B�'b�I/#z5��I��;��� ��K�2lIs�V-�ē�?������?���H
�(�c�@�%��@�h$J�����<9)O��D�O��Ĥ<�2/�-c�)ߕO[\,�V�/<W��`�:D��	��d�I\�I��`�	�QN牧-��i/��X�\h��:z��e��O����O���<��ۜ.�OaZL W�Ӹ(/2��DF�2~��{�'h����'��O���3�~�>��L���Y�ʍF�*y��Ju!��O\��<���13�O���O�`� ��b�F7L6{rϚ�)h�0J�x��'R�-�B|��"�3�_�o`.hkv� C3Vٲ�iq前C����4[�������S����W lڡRn�%%��6L�9���'B�M��y2�|��逘}|��P���� rE�6z��ǝ�>7��O^���O8��g�I۟����DR��
r��p8�J�Mʉ������$�bм�"���/<�p��,�!)�0�m���	ԟ�AsM����|bI���ƭ�f��r��ڝH�ht�`lӒ�LK|���?���n=��+E �0��X�/2�E�iG�M�3N
�O�3ʓ1�`��C�s �l ���,7��mZyyB�'b����	˟��'���C��DB�y�$,@5ީ`�L�>�"O.�d'��?9���%a�tI1W��8R�.J�}4������D�O���O����O^��,�O�7�Ictrl � j�������M+���?�����?���R(��U즭´$Z06t�`��`��;�K��>A��?Q��?Q�t�>y8��i:��']�-�Q�,W�� P�Y��P��.f�j���OB����"\M�,X4�$`ӽHV���(`VT�3�i��'c�'0<u��P>����P��F�m���J9��E�֣W�(�b\bN<���?1�+�;�Ġ�<�O(��y�H0�0��f��"m��l�4�?���6������?����?I���?���5J��m��\������B�F����ڟ�����.�6b�b?]	��N.,�-��N �[�Uc�jg�P\�de����������	�?M��������Ъ
N�fEHQ:��b����h���M��7����T�|"�'ᚁ{��͉u�܄�̘�m����3F`����O��DR.pu����i�O��ɫ?��iՉ�rRb	��A��@�y�"W T������O����#KN�Z��׶ZE�̀�@zp.��'�l�x�^�L�'�|bB�5lB����aD�HL��ap��(���\c�Q�E"�|~��'���'F��'�@چ ����H�$�p�ۅh�F7��O����O���h��y�K�5m��5΅�	�@�#�ߞ;�%���|��'a�'���'"���ӟNt����\�4�ė�~<[5�i~���0$�������
�m��7R�<e��^!T%��F�Ͷ��I����I������`�"��l�I@?Q
;�!!��G��4�N٦���p��ڟ��	�^���g..���;L��j�CG�?�l(Iw�W��ѻ�?q��?A��;�0�#��iL��'���O,�48V�N�&Q� bS�E�5�boӨ㟔����u��5f(4f���`޵"���{s����M����?ф���?A��?��r���?�1��ڢ_��H�C��uW��mZ�����v 	�A5�)��7$i�G�*PK`8�U̖�m%�6mH��R���O��D�O��i�Oؒ�<,�վ2�-�T��,w��+e�	<D_��%!�"<�|*�B��5
M s��)c`e� Zѻ��n����ß�)a����ē�?���~�L�:'����3l]�(
���wNף��'&xS�y��'=r�'� 㑕B�� �C��l�8 �Kq�b���$&q8t&���Iɟ0$�֘�G` k�lL�q���u�ܧf��"?����?����d�=�M�vG�
8��y�ʖ�Д���.D�I쟬�IJ�	쟨�	0!"� &��Ҵ�"CI�|!����5�	�x�IƟ|�'q��"��f>	Ŏ��K���P�G�c ��:�x��˓�?�(O����O��d��>���$��'�z26]�"F3eEޕ�wZ��Iǟ��I|y��H�N���'�?��'X�b`�	 ��Sbbؓb�ϐ��F�'���ԟ��I�hB��`�D�Ov��G�مAn��R���-]�|���i���'_�	�}=�h�����D�OP�I�u���yGgՎ{p��X7��.,x]�'���'�Bբ�y��|�۟��H��.$����&a�y���Yǹi(�� 3��hyݴ�?���?9�'Q��i�ɹG�O)�Z !EI�4X<��g~�
���O� �B8O�O.�>�s�ICF��M"�8#;0�,~��8e�����̟,�	�?�"�OvʓR���U-� 2NT}�E��~�q2�i%.�ӟ'��Q�����|�DIk󌋌K�Ҕ��"�pV�i@��'#�7:�����OR��^�
!1 �ݷnJ��Ӧ)G�!5�6�<��_�S�?-��������BC2���B�r6R�(ed̎2�hTP۴�?��hֈ�?���j��ܟ�$������+H�
�̒=�����4��ñR����@�I��(��Jy2I�2?�������z!^����'��8�Ç)�$�O����O��<��ʌR�� ��l-I��|��H��|b�x�Iӟ$�Iҟ��ɦo�U��R���
�p���s��}����4��d�O��Or�D�O��A��ù4x��Kʤ[�L����"@=��;�o\����O,�D�O��q��3���V���h妃��#P�EtZ7m�O��O��D�O�T�Q�V�6y�h�
�OC Ћ��v��6�'��Y��U�T!��'�?a��>y�9�aEj��q-;t��A�xR�'���!�Op��68��b�IŶL��e*�Ù;��0��>��	��Eh4�����}��yڬ�	@��G�6�2�f��y�*��3��QxRA��&A<�k7C4F�jmICJY�.T��RE��x�+ӝ"���H#Ò�2il)+�D:Z���
� @�K���4ϰbf!yà�#c�K�^�@�!0��%l�Qq��	;82�Ԋ��� �"�#m�� �¦̪E�
�H��I�_9$�2��u�4�1�Ԓy�T�vDN& _�\���O����O����ź��?q��D����S���O����d�SM?�4�Snx���GPH��|)���n��a��C�%�O0����PD�!����{�ƹ�p�O~��@�'�b�|"�'�^� G���w�TLjRϚ�8q�$�:D��0�, �Rx��LW�v���h�cT��HO�Sjy�)�H;�6P�`ˈ�8@��K<��H�;��D�Ob��O\�+���O��$z>��a������7�:4&� Yj\7�����ط4.
("���Kx��ɐ�ַ԰#q@�k*
 �K�",(ԨP�B�9#�U�5d�Xx�ظP��O����	qfvE�� �m"����#�O����O���#d�,��i�$��#���|����_Q��c���7[V���'g�7'&�̓)���ry� �JQ�7��<�(�F99��
�..&9���L/�a�T�JND��$�O��$�~�f��uaųJ�S��/��'Ӛ,�U	��w�����̖�(O@�h�)��D���)˿� �x�Ĥ��m�(Q<.�J��R�D]b� U�~p�75SH��!�1h�NC�	�\��g+�y���#�M���D�`��3k@�T�E������'e��E��牄%q<��4�?����iV�M�Z���O^����V�R1ӹ&O����޵�(h���O2c��g�'�d}If��W��9���T�9����%��R��"~�I97��p*�C@�$��O��K�(�P�<E��'c6|�!CÌeWu
ċ6|�����ʆ� ����%�	,�n�Exr�+�S����C�*aE�6���KG�3���'
�y2�0:��'#��'7�ם�杩Hx�Jd*�@�a
uHB�N�!��g��`$�ؽc����(�?#>� �'��FN)v�sGł��?���8^�(S��G8��3ړ���i���Zo"X����J ��~�(���d���2b�ŷji"	`�$��4�4ȘCi1D��iTK�(:�j���-��*�� �HO>q!�Mӧ�#*m��	s�2|ހ�`�%D7�?q���?A��4\ϧ�?ɚO�Bh�3�5J,\���\;mhhyz���@Nt:b��;[����'��1���l�T1�q�ٵ =�qS�E�ٻ�ē-F@�z��'��#��?	�!�72�L ��Ώ��T0��?)������O��rw�!E���}Db2$MpSxI�ȓH����.���y�g�� �4Lϓ6�	lyrU�&o.6��O��ĭ|�.�پu�w�%�x�S
A1+�H���?Y�M�Τ���\�3��A��"�>�O�B�d!K�iW�M�g
BGl$3��$�)e�B��GO6X��}wK?x�A�����Đ�'M�#��h��Y�6U/`̩����D�"O|�B�-��M_��@k�9Y۸A+��'0O�٘4�ٔT��͛�+A�f�6�#�4O8D�K���1���̗OT�a�E�'�"�'��͐��U|�n�k�)G�\�d b���H��Q��T>#<!㥑��@��-�:U�0Ae�2����G�X�S��?9W�X�~O�4+���*�����͉s�p���?Y�O����O2���-E9~���@�%�佐�>Ox��%�O��@
�Q�p�ÏG�bΪ���ቪ�HO��HF���ǃ�i;�L3����l-��	؟8��À�QP����͟���ǟH;^w���',�9�0"�/M�%P����o:Z]0�'�p�xqm�:kra{� \��@�C:D
�;��Z��~2nR'	�4!*�'$��7�E�Up��S�#Z�Ѕ:��'�\Pq�'q����,O���<I5�S��V��*�9'B�"���]�<�׼>C̛��C^TY���ք����'��$�1^{��m��H�ځ��dI69H����{�,���˟��	՟��c>����|��L��$�d	T>������Ưt^`t����&�2p���K$��<��E>8��Ȑ�m"oIVX`gNکRP�-@B� 3R���b�\��$���O&�ğ'�~���!�1Ac����d�O���?��ʟ>h���yE4�q��� ��X��"O�q��B�~Խp�F�
���5O��'Q�'�\#}:3@W� �@���F�E�!P�/�~�<q3�L A�j0�Dɜ*7�N��ɕ{�<� ̜�E�ZAr#�
7򙻅��p�<�I�v|���6l�?�<3wb�<��dحC���ktW� �����E�<� ��s4�P�y���#vk� Ծ���"Oj� b� o	��I*Ԙv�,�k�"O��diĪ4�ThSGA�o��=@W"OD�#"+��]J�����2�"O`򥏌����,A�BZF�t"Ox(�����p�P0G�<��"O� ��L�e�jAq'�H1sC*��"O�U�N��MV�A���o/���"O� Z�JՓ �\A�,^�mC$"O�i)q�/d[*��F��$�Lݹ"O� !�A�x�����&E�9e"OF�!�A�1�D�/��و�"O�A�gOr��HE,��%�v���"O�A'���9��խq�� �"O�|���̑M��+� {�
lr�"O�X'��@�ごs}����"O���
�q?��	c�#�Y"O|I;�GO�F�q�����"�m�"O�)�)Ӻ#�Dq�f�O�հ�"O޽����L�{ �3(w
�h�"O.�I��o��9H5!H�Q���k""Ovŉe,Y�WI��c�f'V��ɴ"O*�!���|�Ը��dR'q�AH'�'������&n%�!����2@`���!�ѱs�m�R�'z�, �'�NU����:P
qӱ'��_D}���ɋN
D���[*:�Er�c����$�j;&=���S-d=�%d�yKޭh��� ӦT=-H��)�y2@+v�Z��T��Y"A"C΍(��"׮DM�H��OlɓR���ΉP1)YSOP�8fȆijy��(U��3��'H ȱY�_ת��(��Ũ��ҡ\ې��q�[�:��(�ь�>�0<q��\�M�6�r��E�6�r�W����>���9#A�q��U4Y�"=!c��q3��2�eN:3�N���cfY�a&ۼ4�b���d�i��|��I�N�z��1L���O�홥去k"�ơEs����lٜ]R�au ��g�fi�F��F�����T��Hqa%�C��=)2C�J�'�.��a
��1���S!%�T!��'�D����N�8X��� ��2�J�89��Ы��"}���xnpl���{�� �C�M�3�L ���&-����'"x��y�#@�&2F�1�ȁw�ԁ3��A�t��k&k�1]C��ǰ<���e��)1��K�r���1�ғ�p?���FR�eiP!��b�r��H6f7�,M]vx���K���ҨR*m���`��(�
\�v�V�V#?Is�M%� D�S肖+����"�֦�"�D�0h�t�
q�J�m�h�'�!��V�	;:z�:d��9�4��h	gj4�Df�dZ�bw�_�;<�AQ�R� ��*�+|�ƫ4%�4�@n�py��>}B�K�@"�E���#�����a���ClϷw|�4BDj�?d�㟴sVG_�vh��h�G�\�cc�H#��t(�V���cm���S��}�'v�9*�"Mw/��%�M+S�N0ja/�����s��)��x ���5�k�$�v�����\��mb_�^���C�k.>�>���	.	:ƽӗ�Ε>tT��Q�W�0ᐤk,�Ӻ{�'ս�?�S�|'����f��P�v��K�>*Q��D��G�}"�.$hz�EC�R�,���`j�,δ�G��`��ik�Ofhr����yRGJ9R��\21\�0�$K-�XKsɋi���r�$f���g�֕��M�"���ůo��x%E�;�����$�:xLݸ�O��!ђ|u-��&�
f>|���i;t X��ހ���K%nW�͒��D��v�BI8Х���d�!)X2_q�k3&��C��J�GV3_���O�z��`��杄H9�p4**]�!���x�6-?NF��I�X�4���Q֜,��e[�$�Q��Q�4	:��>aP ]�N�FXq�@��t��h���U·��I:rŒj۠�b�n#O�1���C�l���͚M�v��g��B��m:��F`����*��y�Cˆؠ�i �JM?�7�PA�I6�=�<x�qa�jp̉�Q�R��<�\��ǝ; �Q�']�<y�ui�%*�̈�	A9Qw�IL�p�a�`O�QKҘIVʆ�Cm@�;v���O@%'}���-���7�J�ig	Fw�<���&~�,X�P��2@�"���1hB�A���d@�>�@'c�T�U=&\d�I����5�>H��W?Oz�D��4����?��u�.h���V-k2�#�MF8�L.�)Vep���&L� #>)ϒ�)��8�B0��i#�!���@XH
��ۣu*�Р0� v�>�:����@L�<'�+����G����U�hQ�6��u�F�<���)g��a�N���3���Ӱ._������!N�`w�P>kJh{fM��E�K�C����F���S!����48>���-+�Jiy�nӲ[űO�<(�@ �G����ԫ�\l�ݨ��ɭJ�=*�H�v���	�Xd���D����� $�C�r����Õ:n��Q�F?O�)#���N9L���:�ŉ���%VΠ<��7�4}��͌���A.� h��Wg��D����	��O<�0�b9,��!R�Э� ��>����	�bnt��Ȗ8@y��S�P�p�0��.P�1�a�ȡ���)�
��Be�^���eQ�p٢q�2��>p^�0��Oj���[�!��i���C.a�Q��k��`mL(�gP�aB����igJC]�3��=N�H��K�Ȝk��Y jY�Cþsz���J;��2�X��Е*ѷp�J�{S��.5E��r��&=�&q���Щm��PW̾��{0�ۏNʓ ��q,�uG�֬G�J��"��$H�Ã55P��!�̇�r�t�=O8QP�)B,F��*����-�$��5��mK��ؠ`	0y2��A4p��q'���P4;�P��LZ�M��$�)I�e@1�d��"p�*�艗j��R��Qs�	B�Z�b�}��T�'�s%�ԡ�Rߟ��샫N��%RbJT� J�%eL5qA.�� �J�<	d��1�FuP���.J>$QdFL�`�J�s�-��aX�t�v`����"'�!��Gn�$I�cx�J,p�" �X��-��i�OQ>�Ҳ�_�IL9ڵFY���X�,M{ld��`��y�DY��%����b�#<�,��'$� X�n�P���7uϤ5	E��Um�	�a0pQ�DJ���	M��?�"或b)�D��h�$i3ʅ!���iE�`�)��CZ�Vc��VlC�Q�e
@B����'k2Χ^m44i$l��nY,$��� �`��	ӓV��`H�R�k��A�t�<E��ʄRm,��f���J��K�a��㞤��=�&�hgIE�pk0a���f��y�q��p�ؕj�� `I#�I%\����%ƋH��j�a�S�s��M��E�S
"\jASaD��H�b�z3��y�n U��H�� F�w��zP��O,�$��1RД���@�OٞM���ʞ`b�"IL�,�ɤz,�
 ��P����H�"Y�L��'}t�3Ռ��w���Fކx�
��OGM��{�{c����ol��eȫ~�H��9���0��I�����1;���ʧ]d��n�"�&�X�b�$j<M)
ߓn�L���ل]䈢竘'g��k�g�$o�Rq
�eX�_>�xp��Q�S���	^^���ې4?�d��]�
̫ņhNpy����+@Q��Fe��}��̦OV�y��6;�����ɪd �]�&��,N*X�Dkp��HH�5/�zP�欒�4����9�|,i ���6d���!,E����� �Zh&��a�ς&`h�iA2E�+_BR�;������� 26`����k�91��$��lp!a�/�O�ep��ţ[Ԗ(�VN/a���!�'�Z=�Ae��/����PB�dr�{*�rD�!�MJ��� �	�,�507�6D�dJ���+�>�C��X�n��<��*E�D�Lp��T>}҃ƕ�j]z({��E�<a�gĄ�j�c�Z������ix�����	6�FM�cf��r�����Wo��T��<�!מ!�Xyx�͟E���gno�'�ĽH�(�::�}A@NCD�P|R��D1��8�3��.9��є�	T�$
�d򸉔OK+W�x�B`�W��Q;E.��ya~2⑳u����3N(5�h�%�ˏ�?Y�A�?zcĀpUK����j6�S�S��n�L,r%
�&@�|�	�U��!��&4C�)	A"U�F+$�� �K�l@7��и��T�@VI&�n.牂m�����@�tX.��")P#D2��$@.c�2)�� Z�G�E��>]�"tqJ�t%�I�p���ё#R7w ��BS�@�+">1�R��p9#
O�5�,ɲ�z�'h@���{�Ή��R-e˲-��'y�ä �>0�(г�S(�h�:��L����k�<�pL>�|:�wԌ�sn����ᒭ�y��A���g�ص�>nY
���g/�ԍ�=�O����MjV&��e�o�pI�a�|�'BpH�e�'���b]>�&%���S�D�I�r<�  	�_]ܭ�W�	z�Je�=�O.�z�I2n?��Ys�'�D�RAr�����Z+B�h�ETj��ށj�|J?!#�${޹����t%�����3�P�,���)%吖o���J�� )\p�EMPZ��y�˛�mj~�I!ȋGo:1�ҋ���:0�ҫP<��ۢT���O�ɕ~�:��fVE�\���%�6|��x�diC�M���B't�M�Ģؿ+�v���sch�&0���J��9�) �D�I~��F��0���&	�2��5�	����� �x�Fx3r,�Y��ip�ހ�@!�b��?����Fw��3?�e\/lo>��g�+?�tx��ͻ��<1��_5���t��Y}R�S�@�\e#�u�F0Rq ��OE:�
�P�P[�bU�PӧuO�H��wP�ٸ�Sb>��	P:J^�xH>��Aր%:�%?�)�4�!�Z[@2t�@�# F԰LI�&w�0 A��r����C)�U�"��i�8��gɫ��8�rjX�e��ذF��=p�O���"'��-{�h;�N)��'���@7-id���
�!w�:�"B��2���7H�)��1��y� Q <��݂g�/���s&#'�7��(���gۏ{�r0p�(!��>��2\Պ� �K��x��E3��`*�O��Hp��> ��@'s�N퉃�D3K��]�D�Z��B��~rb_|rfH�=?����EP���T���f<qb@��n��J��I% �������'"�L(h�W�DыG���~��Ġa&�
4Ѧ����V�RU��	�pV��2���76�-��sqCˑF��EXR�=.�f��W��k dO�e����fc&O� :�3u�1U����uA�+Y�ՙ��[��1��S�u�~����C�1&n\{���zT���[Y��	��ƕw���(G������z睑)�.�p��n7����W��I����c���16mb�-a@�8D���'H�7|����,�,cD���/��$ٰ,\�D(���T>k���'yA�@*O0y�h'�l�6-	�/ $N$�O�%�����h���8�����'�$%��V����CM�z��ŐS���5I�L�"�w��m �/��`��iX�,ߔj2.�s���&p|�y��9L@�!h�6O��!G�����D�k��CG�%W��Ua� �1O�u!���,[}Ԃ��Z>�p�4Ŏ"��B㉡yĤ�����vZ����9"�CD�/,�\-b#�5��?����=P�"�ݥhG��a�_s<�;τ�U�����S�V �w!�1p%�!Ł�8�n��$�BNa�d �{r��p�2(��	N�p�sC��d�,�X�낮$0���C�
4 �YEx��kHdXⵢ�%�`�I��'����3������+�ͨ�i�4��8bڹ���V���Z����2�H��7���
,F�k�抮kd�#���>>cx٩�jD�&��B�d4�K!"�3ѭ�X�|cdχ�xO�C�	�lJ��(�.�'Q��WeR�=�tqˢ,��o}m��9�&���'i��>Ѣ3�*����aT���r#�6(��*��'q��C5-G�B����B��(����(�ӥ��K�aΓB[z��K>!�(Kn�OlU9�F3IAx��.;)�PZ���:
��٨v�&��0@�M(6��'j,�ve�35��i��A�P�ȓa��5%n�Rıc��H�F�M�b��)$Mv{@�R%������Y-,�V�;�;q�d%j���yR���1���*����Ł�nϫ���F�|~��z�%��<)eM:I����_�zLq��cDwX����֪*-��3h�	)�����ėڀ��@�.�C≩6>���͏2+���{���]l�"=a��E#_��bO�W�'N��Ѳ��`�͓��B�{��t�ȓ8 �SAc\#Uv�X�k���IQ���oȣQ��S�O�\D�r��3XܝbreƩo��L*�"O,M���ΤXfQ��%�qΠ%�����J,J�a
˓�00"skǰ+���Q�1�~���#.��:�j��|�*�(�U�r�^��ȓE�8��4|n��h�L.=f u�ȓ$�.��`�B8:���'F߬`_�}�ȓe�`A���P��H�Cf{�؅ȓ|���#:��Wl�*��a�ȓ��h���K�b`*I�C�5:*�`�ȓ5�����]�r�U�B������ȓ>�6Հ�&ژ�RA�����ơ��U;4e�7L_:��J+�Τ��Ц���!Jky,I�[�O2a�ȓ��`��偟�4�OܠQ�M�ȓf� 5��\&qx�PS�ɦ.�1�ȓt�n-����+�dq� &QLP���ȓC"��z��_�Jf���1I�!�ȓj~귊�<	
tBQ�M<���@+���6��}<�XU��� "O mb�$	bRa�Y�$KX���"Ox�摤+R��a�	�5);(�;�"O�ј�j�\p�l�R���%(���"O:�[k�+@�� q ȁ1||:�d"O�ES���*h�L�b)��0"�H�<�B��#�(��(�?%lmYĢ�B�<�V��:v� ;���x+���"|�<a�@���8����`0lՋ��x�<��_1Q��b��a���A�j�<aA�ʄAY�	�R�ĵ
���&�h�<��b1ιB�04,��z a�<�vo/'��c�&\q����e�<�� �!"i�Lq�K#?m=I���_�<�E�B(9���
X�G� (� '_�<��0!���i��w"\�8gb�T�<��P��c�E ��|򒤆X�<� �i��F�P�$<8T@1}-�g"O���@̅9@��\cIB�=La��"O��{�k>(#@�"��8�09v"O2ei���"<K��� �#��"ObA)3�@#^b�X�u�,$A� "O��(r]�64&��bӡ�\�"O"�HUoӀ���o�FE��"O��A-�N8�IE�Z��r2"Oȡm���`����&�vd��"OR�{â\ hN6��r�*z�*Y�#"O�AQ�_-V�6��%��$��Hj�"O��
�&��J����D��u|,�!"Ob�j�#��� qA�"�����"O0=˕lN9Eg�����$B�X\��"O��w�T.F�l�a"�!��'"OF5��K!b�$D
"�	5����"O�{��W�Go@��1�OE� ��"OjP����
S�"��"X4/Bx9�"O�\ʇE] C������`(�Z$"O��j��O� �g�=$�*�"OHŪ�m�~�dɹ���(<�"O�(X� ΍_�yb �_eV��"Ol�Sv/ކL���u��g�����"Oj����T�X�*xY4ʂ�H����Q"O8i�3�J�
v�	E�M�v<���"O�\Q��^	t� ��F�-,u~QA�"O��1��J���|��
AW����"O`9+���<�0���ߒYڄ�7"O&D�V T�n����K�R�J�"O��rr�U�v^A�U�n�<�1g"O�iF��e�~}`ԬJ.~xL��"O�I�.��!lT�!��$[f�4�"O�i�eh�1E�T��ê»Yd�H�"OT�P����D�H�C�� G�<�R"O6ݡ�<MF��lɒCA��k�"OD�#�r~���k�;1��S"Ou����tX �v)\-,B����"O��A׉!a���HU�<Pu��"O��ad�b� �p苑~+q�w"O�%5*=R��1%
&-�4ɲ"O�i"��/8����D�+�l�k�"O�Ać��B���� շ�n �"O|9AT�U�	�D��I�Fm����"O��j��-ǚP&�#Yx�"O�)�� *W�����DG�N,q{d"O��VL���AYd㚥t=P��"O(�s�fI5J�֘!��Kt��'�Q� �g+�o`:l�ǮQ�n�Q d8D�0A�ȗ@V(#3"��2���"D��!Aɇ�^�X����S�<�
s*?D�X�fg�o:��T��Blz�֏2D��@�IMA\�0��,v����:D��@��]�5��� ��"*wxT���|�#ғ��'����(ԔNtPШ��k܎�C�'�D�Q�Z�	:�`���^�^���'�&130I��<���H�Gƃj�Te�
�'Z�e���5lŰ0��]��X
��hOVв�Q���z���&-�
��V�xb�)��9<\�C�Ɯ�\��`0h�&C��%e�h�tO2�d8 �K�+.TC䉷"4���0��#�&��=��d0�ɓLSb���S�`3��Q�agXB�I�Ef�8�Z�Cu���R/ C�I�jyb��!I�}��ö�P�Q�C�)� 6\�d��l5#wD�g�hL��"O�3ԥ��6�T��ń�#tm�L�"O�MP�NU�5yT���=Q\N!�V"O$�@�CRRA��a�0!��6"O0P��O$F�<A#�ДR����"O���
�D�>=��O�!@�T�"O|2t)�V� \�Q�ѱ"O���1��@Mp�&�ɄD�*A��"O����aK�w"9�S���9�h�R�"O@��mG6}׊M�A��Fg�8�"O���3![>��([�.��E�"ODq�d�ː7�n��Ԧ@��T��"O^�JTGؑ
Yf�@�hX��"Op%9SIK��3��Տ	Z�� "O���6lQq�fQ@��� 	���"O�P�S�HN���[�O h0s�"O��'���q="ͱ"�՗6�:�a"O4%3F��4G���J&� ܖ����<�S��y�Mɝ4��٫��/'��"&�];�y�ʕ�X|9����"%z��T@�:�y
�I�ި�GG�w����y"�AE)��K���I
P�sə��y2ȧ'!�e��( R���nK/�y"`��E,1a"�.]� z&aІ�y2f�1Z��BTh��RqHh�yBlP,
����EtS�pX���y2l�n���1E�.7����J���yb���O��x[�)��8˲���G��yr��`BJJX��q�舡	<�4�
�':�Q�P�d[\��G�ٹ{/��	�'�t<��L:<�lAi���l��+	�'��)����vi�A 2f2b@��'%Ȍ�F�P�@��h�3jh���'��h��C-}"⍛�i�?��kc"O,��aѣ!�^x"U�T�)��%�"O(����8k��+s%�[�p�pW"O������0 *x���N�F�P}��"O��	b
D5VѺ���S/���9�"O��q�K>F�`� R/\��hT�s�x��)�S$c�&���b����q�K�r�>C�I�	���A18fm�U�lC��?F��hE#S _@�u�H6cv�B�IQ[���b�Z�0}x!���Q��B�	=q�	r�2-\ Mb7/�yc�B��
�@Zr��#�&�Jć��L��C�I+/�,t��Ė�Y�b���օLV�C䉬 �0 ���`�
�K��v:�C�I:�Cc�^�+/���Q���; ~C�ɑQD������ zf�ȣDiDC�	��2���	22�RԣA�a<C�Ɋ9�,P�U*)�J��D/[�C�	�2y6iQ�D�0qHd��
C2��B��L�:@�����,ThT��'D��c`LD�mф�K@N�'=h� �'D�d3�W�o���i��8̒D�'D��V�'w��<�׌%u��P�.;D�H�C�:$�&X*cE�I<��óE9D����:h�9�b��H*�i6D�\�5�Z� 4��D�6q�0l��/D��a���:�`��k��M��b��/D��y�(߃Dȼ�Ȟ�FD���*D�(� �Ƕu��=Ƌ��z���`,)D����`jЄ�g C�|���cG&D���A�ptd��S���/֔���"D�� :5@!��JeV���ű \��S�"O8YU���9�`�$�d"O��*�b[<V4�y��9-�僄"O��{c�� O�$K���:���IS"OQ+�I8T�׆��=�©)�"O@�0��N�vh�ɳ�E2{��]q�"O��P�4B(�b��54�|�z"O|e�r�!v�EɅ�$�`�x�"O�0�5`�- ���@�+>�"O��ܙ]|�x��EZ;�N�
#"O�U#��nŜHB�ƈ?� �"O� r_��(|"®�a�����"O���&N{��Xb�E:T��L{b"O�hSs�R(vZLAVC�]�t�
�"O���%C�/�D�����2+Ǣ��e"Op�s�	!?���v�5w�"��3"Oz�CAH�uͼ�����<N��"Opiyt"�\��A�>r��"O����і0���V[=(E�"OZXs�e�э/U�:��U�<a����`0!$E�(;*t����Q�<��M���e�&�l�[/�L�<���[�KMH�T	ʉ��-��nCG�<�'D�/��U�
S�<1x���aGW�<yf��, ��H�" �T$�|�<�vk��6���ʐ�@�4SEP}�<�C��	��)ڷ�Q,
�3�u�<a�J8��
���*M����p�<a�mǡ��i�ĕ�``�I��ih<�G�H#�)��	����S�ȇ�y�.��2Y�E#�)�|�ى3!A4�yBC�H4
��U+s���"lس�ybь1���rCO�d���+�N��yr9Y��0 /MW��Ige8�y��R+d�;��UZ��O;�y� �����C]׸H�
�y��^w64aƈ�f[�����yR�¸KƠ�R��Y��JA�_�y� #.�	`�o�P��AHV�O�y�Q�|���j�Iގ��aZ��yb끼�hcq'W�R��졑LX6�y"`V�W�`lKU�+S)yvBHxV4D�ʵ�3(5& S�%�fP3"3D����Ȁ T��2Mt�<�x#O,D�di�+�2ː�qg�/xD�%D��:So�6��m	U�#�\y�`"D��k���<"
��Ǒv�VhrfC"D�̸��L#~� �^7z�),D�D���\
`�\�p�HݱJ�2���(D�tJ@%��*ޔ���[���%(D�X�5lE�vj֊� ��ٰ�C)D��
bc�5��0�X�J̡ç�!D�L� ��9`�h(��&��507�=D�8+ԂѶ4��ua"��jB�`�?D�+��Ĵ��UM����Э[5C�	_kZ� �/иk��:e�9>B�I�45����F�?�L-"'���@,>B��8)!>,����
��Iw]�p�\B�	�v� �xW�F��@�%�0NXFB�	Ac`:��+W7ldJ��:>�2B�I
[0Ɋ�"�1U�VX"�N�,~J4C�ɱb1B�Q�.ץ]�f<�G�`JB�ɬ&�P]%g��I�Txhw��)�ZC�	O�PJTC�9]5L��M�&cvC�)� Nz�I��r6�iA[�p`�0"Ov�ZS�ЇH����f!�;Nr*q�S"O\�s�Z.�$�憑37t���"O��"��\c�^����_2�AJ�"O���e��rL�3/:(��A"O�(�6@	�<���3!cC�z�H�B"OL4���Z+�&����B�%"�w"O��k�dJ�Z����A�'q"�)�"O*P� ��7L|u��I���"Oސ��E��?����ac��F�|�<I0���f��ܙ6�էm�z|+g ^n�<��:g��S�,[�&�9����h�<)�ꄼ^,MsF$��3N�z��I�<�塖CSB�J��&~,�����l�<�a��(
j����r������GO�<	��ʠ<�@�f��.��1��f�J�<�ӈH6)ZH!���5h��r�p�<�a�>�.�Q���1?�e��Wn�<	W�؋>�9��+�[�\�2wn�^�<i��/B|-2�͚i��=�3'e�<�`�Q�9A^�[�j�A�^,"q�l�<��T�	 H[gS�4ri�r�<����,�8��A(H�S3fL��Yj�<�3`ό2��V�*�Z!)�R$">C��69��qĭ�!z)���W	�
[�ZB�+)�JI��٤H�F�:�����*B�	)�H�K�&	f@���M"t/�C�I�r�FlC&0�6��MK'&�C䉵{�9 a�&tq�%�E
�"qk�C��#eѬ��`��n��	�u��@�ZC�		]d9�v�Ԗu<��Y��J�B�6-���i�e�(��툥 H<x�C�	n���*���Is�M(7  "�B�IZ}� ��T�p�p��2�~B�	+�^5�q!E�
>8y�d�ƨ.C��6_�r�jd�۔L&y��J
<�
C�)	�؈S��^7IAcf�H��B�I2E�l��Ңwm��G㒮	V�C��
p]�����#�BHҠ!��C䉚ja��aW�m ����nN�S\B�I�0�``�'��J�rɘ@Ό�L�<B�I,) �`�#Q�Na��o�]
B�	�Z�ՠ�F�o��Ҍ�0'��C�	�"g$ęi������C�Ɇ�\�z�3F�~�C�E�Q��C�I2��� \'&Ъ��s�O��"OȃCN�Q��%z��sx5��"OpUyQ����~80��'�lE�"O�UiW`͜,z[��8Xh�84"O.��O; ����R�f � 	�"O>-�2-�x��8f	ݬ_��+e"OdY%iQ�Oi�}X��D�@8��"O6ĊT$�+
�^�Y���5S��'"O4N֢>4r�1��OEH�H�"O>�0a@-X�T�2�O�;�ͨ�� D�d8uI:H"�9ip�	�Р��e?D�<�#m˸�Ȉ�$��)��5R��2D�$�4��9�L��Űf�2h��4D�ty5��0+���`�A�h� ���0D��Ձ�C��y���	F��zUF-D���]�/X�eL��a��0�Vm)D�����*O��qZCb��ocf��')D����m�@���Ue۳,fbi�#,D�X�����t�4�
6�ґ�Uʈ4iE!�� z�t��Z0�/���7"O�+�����ı���V��b"OĉqF�%�N`�5�jɮ��Q"OH�R �OJ�dR#$�:1ɬ��!"O�u�H$v�f%�։Ɍ+�u��"O�Y8T�E�;aꄢ�j�	Y�DL��"O���X`�æ$��ru�M�U"O���H�W�D)�-�(cIL��"O�52'ʲe~f�S�L��8"OTe9�nO|M��d�5Ϣ���"O�PcuHQ&����ׯ�D�ܴ��"O�8������e��3�"O���-W�2��t��C2,�0�!�"O�5h��=�0���h�H�1`"OJ�k#��'T��P��8/и��"O����`F�=x%�'�3���"O� ��!��.��E��?B��-H�"O�ذ3)]�{��y��cW�.i0���"O�p����ֈ���4<NJM�"O����Y�p��८C�h��|9�"O�L됏ѐ`�B���ũP�>i�F"O�b@U���9��P�T쬺F"O6� ����^��)����%a� =��"O���(yZ��8$�ē8�d@і"O�4�@@ɸA����d��I�t�C�"OF�J �=*���w�S]�J���"O���4D4�����<A��tp5"OzL�f�+����� �+��""O�\ˢ)̉Jk��'�L �*��"OTEQ���g�=��c\�]�dI��"O�\���Ȟcb���A�K �x\b�"O�|��ϊWg�	q� B���P�"OP��.ӭ
J
��g�& �za�!"OVY���*aY���r�h(:""O�k��ڂb�,-�3��l%J)��'�RPcp.)7bɔ�͇}0�C�'�A!��/V��=rg�_ JhМ��'������ 5J����VI���q�'
L�����?���JFӑ��r	�'���j��!y�z��������'jԨFb��lA���Ph}���'�����Vp�x��fϦũ
�'�tz�M$���a�ć=`���	�'>^����\�f˸�y�G��_⾡�	�'� ��
��EB(�Ia�?K����'�ʌ nޠ�02��ۮEŀs�'T�=�1J��fU���R��'<7^�x�'�P�0F��: ��Y�
�2��'|�S��\t�@YE�*{����'�lPS��zV�e;R)#��5�'�j\Ȃ��:4�ui�*���i�
�'��*U	�\�3�b���	�'ϊY���TW�����y:t��'�j�s6�Wm șR�@T����	�'�F���lĮa8آ�K-�Z$��':$�Z7��r�P�eшq�dJ�'vR���Ono���5�˲k� ��'��	��f)3���$΁�N^����'�~D�F�Y�Y���C�4mJ�'rZTa@F�;!�(1�Ĭ�%>$�:�'������̻"����I+�J�'1��%(�$��Qq��˃D�4iQ�'�Q�RY�P@�I �:��T@�'�8� b�`��d��Ҩ2J�4	��� ���&��fT����Ϫ1T*��ȓ͐yr�BF2~�3��D�	�D݇�X"C�d$J�2�2�˫nKX��9}$�C�7tY�|J��]+5��͇ȓsĆ��E����(���ͪl?����P��4�5Q�
���.e���ȓD�2�I��	�T�$���W�Xh��k�Th�e.��&�t��0J�͌m�ȓl�0j�ʊ42��փ��),�l��@]
�r 
	6�:��ˆ�}��9��)��X���D3 X��u�N�,��ȓ�F�:sh�Mi|u��F�z6(��LO6��ũ��0�=��B�֞���(-2!�g�RJ)��bFKù]��x��s�|L{�=Ub=2��7J��A��c��@R!J�躍`�>�
�������aǯx�.-���ϲ0G�5�ȓj�(����K�Q� 8�̠�ȓkQ!�ˏ��J�RE�A�p���ȓY�*�DL�	��8�W�j t}��S��	�F#��
3T���&ư#��ȓDj�	�\7'ʄ(2�V��jt�ȓwd&aX�O�vE��O7eϐ܄�g��tҡK7-]68�	S.SY�e��
����?k�1�5�	nRՄȓ<�(�s���!!C8u%��L?��ȓ�6����ʹ��Tvm��^����ȓ%$p�����2("ԑ��$[ �n��ȓ>u��"lD�I.Mb�j�i�ńȓI��E{�A��Y���QAҬK:��ȓ!$�I;�7�A����g�U�ȓ�(C@*�;w˰8)t��_8��_ 	�w턕Y�t�h�+�L���R��c�	pg�p��lǫT����ȓ`$`��)�t�2у��-scr�ȓV�F��Q-ԤӄA5��L�� ג))4@��?�����ۓ��1�ȓG�ƅsGJ���*��S�1��H�ȓQ<(d���ƿ���ɑ�4��B�I���y�-���[�B�9�C�	�Yx��jT��67����A$�:M��C�I��d*�l͡\�Ҍ
V�=J��C䉲n(�ۦ�^9���*���4N�C�+\Fv��VK�(}�z�ز�ǌ#�B䉕j�¡	%�2-D�)Bb��Qݡ�$5��5B!��Ct�m2��Q�7!�$�';I�d��.'R�p�$l�
 $!�ā�:(~�!QN�lƈ�H���!��1�(\���!\�n���7S	!��hx�����(]B��-�:5�!��l����&͆�kx��u-��y�!�dF�]�<���Ț�MFv6N�=C�6B�=#V`%%�$�9`#n-�B䉚e��`a���v��4*d����C��	���tBŕ@��JT-V�aj�C�	�p����2Cך��V#��C�I�7�|0��m��r6h8`�S�MP�B�I>TD���'�/�d ���XB䉺"�Z5�� W36~����X�k�4B䉷a�BXa��}���E�bg~�i��"D�� ��&�l�v�w*@K'"D��Kd�%>ְ@W��p0���2D�$C7�R<�bT�@C�x��qS+D�TѶ�4'�����r�L��G/D�� ��:3,L�l�~� c�1���0"O2 !�Nt��
A��.����"O@�#�]���I3�]�!�T��"O�쓀�͇GF\��
�(Q����'�ў"~B�b�'����耕R8Jl�`�K��y2�ݼDR�l!G�0H�tı`.��y҉����h��i@�G�v�`����y"�[� ���P2��7?6� ҄�y�$�od9���ߓ5j�ҕ�5�y2��r=x"GF(�|�Q�ޏ�yb�Э=e�m��ϝ���!�� �y�nL8�eʇ
���z�P��;�yF�2�1e�K����'���y$�; �XuˇOPzŠ��Ūʨ�y"��q.��K��Z0y�V	+�����y2��L!����cRyA^�j�/ȏ�y��R�j��i��d�l���2�yb��*]F K���5]����ǯ�0�y�Њ���*��=P<���`���ybI��m�~A���نM����k��yB+G�lc2ŉ��;����AK��yb�;۰���h-.oTMZVG��y�(;)qL䊅k��16��6�yR*i�H,XPfժX��k҈�!�yb�U>V$Ő�DZ2v~�J�lؼ�y� �W�MtEvd3�E0�y2	3�x���kM�m�J=��HY��yB��~Y����ldT�C֢�yҪ;"f�$[���-`�~�)���/�y�	�%e���R�����Cې�yRh�k��!ɄU`f�PM��PyR�˜1k��H�C'::�����S�<i��̝b�@�*�m[�4Xl�N�<QP,Xghe �\8cU��T%D�<�G
��m�0���K #��@�<�Ǘ0[qx����.l��ړ�R�<��/V.#�^}����$=��@�f�P�<�� �z>e�!���2�( �K�<Y ���d9ށqu ��8�a�E�<a�G��I��1�
�w8��I�.~�<�����s����*� %�R��w-�x�<�r �qK�Ht�
�7�8��"O�<�p&���2�:[ �	��E�<A�,�`~=�s��n�Dȁ��G�<�s��a���F��e]�C4�Tn�<QR�=��P���J4�"!�)^s�<�3�V�z�U@@�ލ*�\|+��o�<ɡ�G8q�<�	�H_�R�9s!I�f�<����k~x��K" �j�:AOG�<��J�<x�����t(8Ĩ���<�A�P�>A��2�J���"��6iOs�<Aҫ�_=ڱ��E-0�l�T$I�<�u�ذ	%�zC-B^p�2�d�N�<	Wḧ.r��NM�ifY���d�<����A��鴅L�?j�����a�<���;Cǔ���O�<�>]���\]�<A�,^*1�1�#۴Ԫ"�s�<���M�D1|�+Wj��R�D����k�<�3j]���i
Cd^,0��t*�'OQ�<�r�H7D���� ��7Ţ-T��g�<a��оeʞz�@
?�8��e�~�<90c�)O�>պ&!��>=֩!W�Wy�<�&e8<��Ղ��ǁ5Dn�pDRr�<9S��PJ�W�]�\�Ka _T�<� �<��Ӝ3�d@�Җ/Hؑ�"O��@e(D�%Hi��D��9pA"OT�u�R2(���u�ۀP"O"�0�@@�_���ѓ��,z��h;�"O�Ayq�X�`-�p��A�=���b"O��լ~p�y#��*z�*t
4"Oj���J���W�\��\�4"O<�
�F���0"�Q"O���G����v�#A��2��D"O�����?x(܂�-T.U5"��"O�� r�hZ<�%V�~�hP�"O�ݩ�ІbF�bF��P,ޑ�"O l(�N�T�P����BJ-i!�K9��M��.
F�Mˡ�' !�Dߓ����R"��"�
��_n�!��]24��}�͹p�:QA��AN!��[��9��˙�A���\>F!�D_�[�@Q��-{f�`r@��$[�!�$R[�~�)��NgML �-��!�H�3v�)�e��.WH��3U�Ⱦm�!�\ o�ش���]Q6���녌Ig!�䗘�x�@ڮx���au!�\�5�	�ʖ�K����q��;u^!�Ė72���B �߫f�f�(b��!�D/C,z|��M_��A�5g:a�!�dK�B��5�F
Dd|ve�t�Y%�!�ć3"�RQ���pj��c΀�}�!���^?Ze��'Rw$���j��J�!�dP>��}�B��k�L��A)�!򤐟|<��IQ���(P�dg�1 `!�d2�&p3�jpD8;A�@?H!��J�w�&u�"f��X���q4!�$�@=\M�p.	#OL\##��8/(!�DŁ7�Px�m�dY��#E��!�$�11ج)����)S�������:�!�$�>:��Y+��E�gA��SD�E�r�!�Dɑ#u��6��)\&M��k�!�D4~�́
���D��G��l1!�Ǔ&�85�6���UAH(���@!�$ZD;��)ʄ�B��d�*!��&jw2�q#�L�J���00.V�U�!���1 ��#�E	yp!X�̙�`8!��F11�<�*�g��l ������m7!�� �={<`K�
�#3�����\z!�D�5KF��A�A�etl
��kp!�D��O�t@�]���E��-2G!�d]5\hPy(1m��$P#'�.!��� =�0U"a	ۚ���"�Ӽ!�mH�%Ѐo����u���4!!�ԩ"�H�˒���CLP*!!�DM,j͖�at�N8:�6MXvi׏n!��W6���
:�00Ti� ��'�ў�>�j4fG$r"��W�@�A�2�;��<D� ��G\Z�����0G��Hq4n?D��Zp*��r�DUv�_�1�v�[֩;D���b'R�	�B��T�	, IY�AC:D��ʱK��}���ܥP��qq�6D�P@X��s�R�n���0�
-,�!��)`���c �~�������!�DP7��kU���DT,#!��@�p8r�H�:4�������!��ҬA�ؙ�ۼɴ�b�E�5<!�$Oh�l��w#�)E�x� ��T?o!�$I1e���e� :�R���1
Z!�� "$��aް�T�����z��@�Q"Or�A�DF{�p{�`I<� �%"O�����H����PS �:>�)a�"O6����.��tB�/�uFr�"O�`�'�ֆSê"D�Q�Y+�0��"Op�*t���+)����&�݈"O�l�ac]�T�$���Gɑ_r��Kv"O^-×*I�q�q01�1\�جc�"O�xH%�)|	�����-���S"O���6��&���	օ>�4��"Ob�����9�$M�w��(���	C"O�Q���\�� <RP'D��v�h�"O0��M�G��Ȳ��l��*�"O�y��$^�ifjy{B�EԘ��"O���`f_�-�p8��GS���G"O�!:�">k{����&ϝr�Fa�""O��J7p��q�c��o�����"OH#@&J-NHH���`@��"O4Hu�@p;�Кtb�C�N	R�"Ob��"C�J�"T��&Ӆ+-���"O�A�v��>D��P�/Q=/@��"O�a#C�Aq�5A�T�4T���"O$yk`R�_J9���$ZS���"O��t�̜.�����<C*Q `"O.C�N>%n �a�}ArIU"OR�R	�3���$NG�(3�:V"Od�Qc��$wѰ��a╺lF���D"OԔ�䤆_ȬxB�� ��0*O��@3�n����F�]��Ld�	�'�j�a�h_�>�3dD��Xհ�'��C���Q=N=r얣P�T�[�'�b	���@v�!�qfY�#N���' ���"D��|S��,+��x�'�(�`��O1jk⇕7ܒxS�'�e �퍊g�(A��͒z���
�'��1�PDS�u,���\<j����'�fI�V&�9L����T����R	�'|�I�R�X6������ux���'5�ٻ#I�*�4��d�hOx!�'�FTZq'S	 n�QT��.d�-�'���!�X�$	�:���C~qa�'�b�Y��Jn�Q��L�=څ�'D�t�"ߴb�\�ـ�EO�`�B�&D��Ӗ�]q����bE:p��,�C)D����A0:�aS�W�n��0�%�&D��c߶%��\��	�8\ʹ�Q�C9D��(����r��dd��_�(�aO7D��b������e�O���1&k!D���4��?U'|��i.cGr58"�?D�`�$��	�M�R�T�r�(�V�<D��˵K¶]"���� t(��d0D���rə!$Zݹe�]XT)%�,D�X��QbaNI�ҋ�a� t��%,D��
�$B>z�"�{�Mh�,���+D���w�
	$RPZc�0����<D��k$��zZtH���)`Ɏ��Ӌ:D����ES�6X��)t�Q0�@x1N8D���#�$HD0� F�SK[���K8D�X	�H m�j�&ζf�4�pUO6D� ��� úlh�"�#� M �6D��R�(��C������d�b�<a��ͭpy&Ƀ��,)�,�`"�[�<�7���z�x�iFO٧h̠h(���}�<����XJ��P���J��Ət�<� l�6���"1���`���R"Op����%���xC&X�9��0�"O~�x@G��Up��HR�A�8%s�"O����I{���ӓ�A�S�.��4"OY��$�	P�Θ3 �@!jfxxц"OX�bc�tɎq�#�V7k��җ"O(H���܀K �	s�'a���F"O��2f��4j���� G=�ʥ�D"Ovɚ�hR5w�^Q� Ǌt�<��"O�rdܹXD����'U��m�"O2lH�ȓ{M�������H��"O��@�E
�E�,��%Ҏ,�Ṳ"O�Ѥ!�>�r�j�#FP���["O�t!���>V1�ؗ�S��j؁"O�h[f��84�|<��V y� �;�"O|�b��̢""�h��?�����"O�UK��H;;mda�
�#�&�җ"O|p��1 ���$<-[S "Ot���^���C���kI�xP"O@,caa�.H���)�Ʊ�8!"O�i�3�_/^-�uj0	Ӱas!"OQ��m��M�d̀�����|���"O���&��)���Y7/��%T"O4�I��X�t�2a����*.Qf\P�"O�1'͜�K�q���*w6��@"O�miBN��.�}b�	; �m"""O�%(v��RҦ�*@Y����y�A�8��0���3���U�B��yR�ؖxj]H!/��)z�0�	���yK�F��(���k̘iE)ǎ�yr�>}w�p��ܓV'�`��X��y�Q,XB���F77��m�ꘀ�y"ȷ7���>+&ޜ��N��y�R�0{��rS�߭3���31l�yB�	�F5ZЪ�)X�WT�| R9�y2���������:��0����y�8,�b`X��;f1��h����y�g�|�܀1�Ō�`8J�I�͒��y�'�#<B
�_��A��-\��y��ՙU怼*T�]��Z`[��V1�y")>����w�ǂj7hPc��F�y҉�=����)�(0}�`�w���yR�T�M����ш��"�6�p���y���B���yT�Z�T�Ц&� �y��kTB����S&�T�J�j�*�y¯�6 _��r�^���yD
���y�ą�:�}�E~�\�d���&B�I1n*Ҡ���$�[#��2>H�C�	1]b�9T
��K�b��M�X��C�I#@B^��Q�� (欨V��6!�XB�	�he>sҨ�	A�P2"�X&.�:B��1{�y���͗Bs�����'��B�I�v$���KȪ>��(�j�"�FC�	�P[��J�t�RT�O�;"0C����(����%<n���Ѻ/9,C�	7o��� b��;5�h0	��T� �C��'^k��Qf�%C�@pj�ɓɰC��34E�A˥$�
�R7��,i��B�I&H�J䈇^�h���I�v]�C�If0����	�Wb$���KϘaBB䉀i�(�*$D�k�L��"�A6)�C��2r^�3G�	��R��!!\�T�B�I=X��D ȑP�t6@�JB�ɝU� �`�ٜ!
�Z���8,�>B�)� �-�R��c�ܪ�n�(+Hp"OZESF͛�O��ZeC�51��"O:(J�G˻?�$��Sh�,|`1@"Or��(C��°�'E�6���3�"O���u��0k��a�CJ��b"O����Ə
Tiz88@�
���"O�4x� �&�*T�`c3f��R@"O:�1G�_�&@�<9��5�%f���y"D\"z�T20*ԟ#N.�Zu (�y�ɉ�\f
�p���!�d��%̞�y��I �@�v�$�v�rVdY��yBD��$����8s�>U�\0�y�j��BLj��e�dW�����!�y"�I�؅ ҭA�b�b���H��y�Ʃ30<�zq.نX�@�u����y���"
�527�W���3%mD?�y���``Kb��H f�Ju+��yr����ư�a'Әu j@{�OƎ�ykx�]�W���Y�CG(X�C�I�h����E�ą�������zC��`��5x$�H�D98���FZ^C�I�5����g]<�y�	�%{$C�	�;��A�� �~��1��;O��B�I�W#t�@���L��&yG�B�(a9QO�-+b�pa#�4#
�B�	+s��QT���L�Ц�LBRC�	�qS@��q��:K��8� Q�Ps\B��/?�X��g�R2t��D
�A*.B�"LW�4�s�ºt�h��B��N�lC��5�(
��[�Xul� Gm�4szC�I*5��jb�LOJ4�ABŻ.BrC�I�$w��afA�0Y4�p�M�/�C�I&v�p�e�O�Jl� ��W�C��:s7Z� 7j�+G�rĒ���B�I�	��ҢL�1V򴙂�o��B�ct���jC�+�����?K��B�Ɇb�ʉB��;0B�����MM�VB�I=^A��HP�L;D)�pƌC�� bH�2�/~�T���_�ZsPC䉪%?&�gK�>p��ʖ�%�B�ɘC�ƕ
�.�.O`t0�TI�;+0.B�IL���a"iWE(4j\�z���"O��{�0L��5[Ý<Z����D"Od����N�OT�N�.���"�"O���M�����#¨j�j$"Of�{6�X�d�xub��}�\8;�"O�XЏ_�EIY2���m���"O�Ī'	B?!7�a@�)W�6E3�"O����@F�IR���r�a��"O��Z�Ns�X���n�{=�Y�"OB=�e��=+��16��?'�s�"O�|"�(�(���1"�${<���G"Od݉Ə0A���&�'2n���"O�S�o|�E���X�L��"OT X�D�2p�x*�<d��"O�,�g�WbPd�Vo*<�5"Ov��s�Ⱦq"��IѲ"O$<��'��	@�hpk�K���Д"O��0��!k�`5k@G�ޜ �"O�Z�ŒZj�hx!�P�a��uC�"O��
Ղ.����jUN���!"Oĝ���lҖ��U��>�zh+1"O���Je,�l��h@�W�29 c"O��X�C�q���!`�
+C�ا"O� HQ`a#�JvI����,� e"O6(���M�<� g�'u�<A�"O�L�0�ڪew���,� =ba"OXt����qv �z��*0N $�q"OJ%���Lm��A �ň0BD�Y��"O�ي�EY�hE�r��d9�e��"Oh��A�ې{�Z@(��/}\]["Oz����8|c`���c��ON��"O�Kr��y=����j��G"ORMPD�K�#���3"�Χ	H"h�@"OPT��	��y*rh�6�X7��8�u"O�]�pa��:�%��0y�%�"O>��4-�(K�`�ʩ^r�eT"O��x�� CjD���� {pt��"O�$L�%����+X���h�"O���@�Y�ZR�]8���s"OP�J��YY�X!���T�Z�!9�"O� �֡�^��Dc���#{-:�x�"O��ien�|��4���3-����"Om�b#�4�ZL�ʕ�w��"OB\p�#�"�+tF�d�屒"O(�*"m��v$��2#&L4q��ڦ"O�	�䘌,J:E%�[��R3"O���!�o5:L��E�~��;D���d�?rD���īC�b 8�&�.D����?��w��,?&*�BvG,D�4�c��3$�(I�.Ҹj��P6(D���0�6�;�!Rg�}C!D��� O�=@��4���̽ �Xy�gO4D�(!�X�O�``W�mh�i,D��z�&\�����v�̴J��;�>D���a�J,QHN9��$&��<0�;D���g��B�$Z1�Et`;T ,D�`8�D�!.{�qdʻJ,�I�<D�8�q-a:8 ���\�KX q#/D�p0��BO�-���ۤ�4)`�D8D��#goJ%;��Yk�,�-Yt��S�3D�����%~�D��vmU�w%5y8!��B�XZ�D!S����"JՊ!���*G��՘׀�0�E���$d!�
�
�cE��1��|�g�A�=!�$�o�ȠG!�Tϸ}�cK0i!��&mǪ�2q��w�,9��C߶!�BC���w��k0cҚdn!�_)��EIBf�,���z&#��D�!��6p�`���.Ә]X
ɻ�`T)n!�DD�6-��ٲ �%=�અ��k!�$���j��6f�)m%�5�c��h[!��R�`4Z�ՃSj����_iN!�_����`䌖]rH�k���:�!�d֯[Z�@�ENpΉ3CB_�ee!�d&ppR���@&QM�q���gT!�d��2Ot��'��2qg(頰�^;h�!���H�t���C<;�P1�F. �B�0g��
C�I��"�C@�btC�	C`�ɚ6P�f�$�R%��atnC�I�d����G��ƅ�(�B�ɊƆ�B���ǜp� �)7 B�I�Zۀ��d�G�r,*TEN;#j�C�	�G��Y��,S){@�H��:��C�I��4��E�>X��h�5'F&m`�C�	'O�!�S%N7G���q��5#��C�	)ov$�9Ĕ�Y����Pm�3O��C�a���H=:a~(b$W_6FC�)� ���f�F�HfpBF��N�+"O����d�;�M�����h��"O���(���FΔ�9R��q"OJ���D�	����/�Q;ث7"O��9s��	V:4ő��$H��V"Oԁ�Woźyഄ[�N��`�aF"O�L��9a������t�+ "O�h8�ā1��T�'ɤc�=[�"OvD�`\k'2���T���0��"OvH�w�Fb��*k?",c�"O�QY�A�Y H5Ʌ�.Ș�ڣ"Oz�zS�ǟ�2A�B�����"OΡ�#��uX.H��&)b��y�"O��p��e��t��oٱcA^���"ODCt�l+�Q{A,��8���c"O���0��3w��5L͢i���ZQ"O ��AE�S�8����W���{b"O ���HN3q�B�֪ګR�.���"OTy����4��g��'�  "O����t��Jf-V1` ��:�"OȘ:tlF�F	 I���)26"Or���K��I8r$�c)Q�Q���S�"OL�@��;"�\(�g���"O�-(b��"|<��u�G�`���"OB�	W�  `�&�
�Z�p"O����e��<qJ	Z�E��N�$1��"OjiK��Ѣp��y��t!�I)�"O���G�R�n�`� cL$��x�"O8�b@�5&,�P��∗3ƪ��C"O�����Cs\ c�P�{�j���"O4a�G�#4�L��E��q��Q"O<ԑ)��U:7���F��t7"O�e��@ϓ/��ȇ!�Mi�]i�"Od���
Y�P�Up�U#. T�p"O� U��l���5.G?FŌ��"O 	!��#^����2�Q/8Ad�p�"O�%Z�*�0�G��S>����"O�萦��uʲA�f$�U%�a�"OZ�3#�>��\j��)+|�@d"OE�a�߽P�z��EI5:nՈ�"O�UzՇ��a%��@G�Ǎt�0�%"O�(!�Hv��qQa圣t�LEb$"O��PP �2X�=3&�ײG�"� �"O�� t#�����ď0�.1�1"O��-�^�@�q楓'5n")""OV��ǁ/n�p���_$bTq�"O�]#ЬJ����[QK��:����"OL�� �B W��x��$5T
Ќ��"O�ia"� R-�u;���yN<��"O����4YN�=�N�YPp�"O��14e�5�L	Bt�]�;��X��"O
�0�Y"J����dZ)�*�@p"O�b�E�x[
��t@����{�"OT��L|�pMA􀑫p���5"O�!���B�pŶ�aD�C 4�Xq"O�)G�e��!iـy2 IK�6D�|���^@�<Q�f��Z,I�p�2D�r�`һ'&� 4	�l*جy�;D��Q� ��^V�z��5Y�Xz��+D�L['+�*)A.y+V��C��X�/(D��T� r|�I$�[r�hJУ%D�zc��:�P�X��)2I�T��$D���nӷ}�½��ϲC4d����#D�h��1Jy�l���KC~@�#��!D�� �[��z�ˡD2a�D`�""Od�RL�	Qt�i���ʊ�j!"O�Ȃd�T�MR�= �̛:��;�"O�Bw��!����ԟ���"O�9wɋ�4_DĚ��C�q�����"O� ��%ӶH�����x)Р"OLQ�nµ-��
$#����h�#"Oj��A+I ��T`�k�&��e��"ODMx�[bΌ��V� 0��9*U"Of]��Ζ'5��=�’�%��f"O��A�͘�$�<�9�Ǟ;b(@{2"OJIɳ@ݗ ���䥐�YDbi�'"O��Ʉ��qs� ⓰>7V�Z�"O������K�+�R�J���6DQ^�<	��˟8\��/Z�U�U(sFRV�<	���-Hx�6�%P��d�c-�Q�<9�[g�$@��ػZwMP�#L�<��hތn�ؠh���a�8\
�\q�<���;�&QCP���:�"*D�<���ӟ[K�H��J�#�d�;#�A�<�d�̟� 9�)K�2d�BgZb�<I%C�R� �,�ˉd?��ȓYx���tg�<(�\�I1jܔ^d�ąȓ>5���j]� D����j�l��-��Qs��$�ӏO���Q$�[�1.�цȓDw2�8��48�����nJ,a8:Q�ȓE�*%ȃ��,eZ�K���q[�T��]�V���F�a�XM9B E�Eg�Ԇ�b���V�?K|
yS��8�H�ȓFlK�A��`�	)C0i�ȓ�Ҭ����[_^(@�/��.�	�ȓ,P0qew�H��@�{)ph��yt(��#S��hXT��ȓ*��Yģ�1�&��� &��͆���[sM9Q��3vcߥ��D�ȓ2�Z�h����*��v�$/(�ą�I� 	�$n�u��B`�؅ȓ^4hP@oߩfGn�t�̛+�хȓYG��c�c�W1��5��lo�ԅ�_CXmb�k�_�� v�؉W�����NZ~�2D�-L�jԚ��;A�!����@�/W6T^�1��K<�XH��M q�B/���҃U�p��Շ�$����T(�Sj�2��1P<)�ȓ_~�ʄ��s��P"�n�8Q��$��ET>p+ڪYh5�43[p ��ȓD�Աӷla���ӶE�.Y�|��a��`�d܈~�����Ò�9���ȓs�0D���W� !�sh�	E��,�ȓF�\�k_�?�fi�2*A�%��B�I<A^j���Ǌt2� �܀k�xC�	��ID�՛4�*%t��(�C��P�p�삎!�`�I��)\
C�I�P&���HۦW^8�2�ф%��B�	$s|��""ڊ1mLd�����{k�B�ɴ}�b=h婖;#;B���.Z8�lB��$~���c��)��bb.�5J�<B�	�U�ተ���w��)2nJ�}�B�-�te��W�J�d ���&s�C�	W����a^�C�n�3�耕 z�B� W� )EiW�u�*S�
_ e��C�	!AQ"���`Z�3�B���*2��C�I�Mm|� �'����]�ŧ+m�C�I�xy^�i��ߧG����ă=QhC�)� �x׉K�T�����P�$�l!P"O|+`_D^��!E�e$UX@"O�0!RM���<0p���H�@-3�"O��/��Ca��V��(B��	��"O��ʁ�Q?z7$4��o�O����D"O�����|���N[�76�\J�"O��W[�F��9+׍Iw�H�"O�a�/�����m�t*�ƍ��y�lBA(�аeY�k�ّ"* �y�+L* �����`:2܈�i_=�y"�0gG������*�j�As��y�ĨcBz���"�������y�� j�����d��M8� X� ˦�y��4��T��A�/KhޅС��6�Py2���9�B�QG��X�xEa��X�<��(�z�*5���x���3+�U�<їNP�Z=�`
Gj�~��,�V�T�<����:=�A�E�'/$i{��KO�<ѵ��#��ӗF����K�e�f�<����8���d�l�Ĭc��k�<	嬇T�p� r*!��K��k�<bc�U �C�*]/u9�xs�f�<�p*�(I�\bs"`px�%`�e�<�Ġ�-ALUs� �^�A��]J�<�N(�-C�h�QX8��L�]�<Y��D	E*|�{��-��u�H�o�<9w�M�~�`hґj	_G��X�]l�<)�JR9f��p2O�5h��H�m�<1�K�t	�eD�h(L�b�<�0$P/(A#�m�79�:	\g�<���NlP��Rs��e���@`�<�2!�>@�����O�.B0��N`�<���X'}D��x&G�%?&l��$_[�<���<z
���V�F	
��b"��X�<���7P���� �r컠H[T�<9�'�m�`����'H�}a��Y�<�
H#AI|�Z�#Q#!�. F�<�!@A�E�@$P����;�|����Wy�<�c�ƌW��Ъ&�3!Np�r�{�<�n-��9Y�fwt�F�Nu�<�Ai `�ޅ�Rg�`�@�ΜF�<���W6����\�z�����Dg�<!��۾p`����&V��U��MJa�<��D��`lՃ�?1�&T���Y�<�ޮv��l�d�#�$1�t!j�<��+�x�~s�m�*�H$�g�<��a�X�u�,/Nd0`�a�<I��7k�i��٨N�x��^�<�Gw�dQ��A�4�JOp�<��䀼B���S�~�X�
��`�<A�Mz�D��Ơ\�j]�%oU_�<)U���(��"`���4΢TB$w�<	��T�@�X0 `��.�u�x�<�@�]}�̸�G�Q̂�TK�<9�O�_�ȱ�(�~,n�a�IJm�<B�R7�ƉA�k�4�X5Iqag�<����;���B���w�"�����I�<��e�(N��;@.( X%Į�]�<Y�,8� ZVÙ�N�����Ā`�<AP���
X���&��0�"ԫ�"�]�<!w��=~v,RB�I$�&�[�]�<y���e�t��ՠ�#Y� �)@�GR�<�3%ԢT��pѰi^!M�JUѲ-�b�<�3ʏ�������^^nHɰGb�<� �e9�ݴ+�F| �+�3 =@��s"O��P4M%L�H%�jh�"Փa"O)��f��@�e	�3M��Z�"O­�E���̬Md���&L�T"O�Y��dI�k n4󁈎��ř"O�a��
Q��lp0R��.G��a"O���O��W�fx*nƋ,�UIE"O�1ʧ%��L��"�L��>����t"O�U�Rj*@H
�JD�I�]���r"O��U�Ef*Б��ͅ^|bX��"O�t� !W1 �bs�Z$[n䈢"O�]� HL�1j��5ɀMU�MB"Ozũ��/~j��h�52NƉk�"O���ܦ#���p�f�PG��t�ȓ)��q�/��>̴�q�L�7:|��Tw��ƨ��{�@��U�F�-,��ȓC������K"$ޤ{��@QM&�ȓP@�Tb'A��WƠ�"$��O�D0���"Ը�Ǝ.nNz�:�J�B���(lt�Gmj �wF�U
Э�ȓ;����th��_䑫 l�:I|���L���RK<z4�ڄ���5����w��[�iU�{��dI'�	�7Ѐ��0UB�&�Z.�e���\��2���G�z񓣎��R����n��/0�ȓ(^L��aJ8/}(��爻Y��͆�bl��H�;_�,���B�dR1��]W,�Qq��!*W����Ԧ2���ȓ�p-��B�e�
�����ny��uk�qp��ʆ-?$19��)q���[�L"+�i��g�#,�"|�ȓ<W5�MЪ]=�es#K�!Fz�D�ȓ;�0d��eF")9K��P�hh��z;D `B_�+4�ٚ���@��̄ȓ#����WeNA�:�� lM)IG����	�<�yrn�(YM��Ɇ�"�R���GTh<�B���8����n�F����	�:t���K� Y����H$j�蹅ȓa�����Վ}�6$�do  Xx��ȓ1#������A�}�CUa�ȇ�]J:pQ�]y�� 
�#��ʒ��ȓT(����&M7^@Q�b�X�������v����	��j��x+w�^�<�4�,}8J �L(t�隀e�r�<Q�'^�<���P`�@�$YC���S�<�e�#[Α���.0Y|kSj�e�<���N�a� iT�P��p��Ne�<!qE�AȌ��D�22�pۢʞb�<�gD�4}Ό3��((��%�X�'�E�T�X'WQ����Q�H����.�yr\����t�R�B�Т��N�PxB�i�8xKU� c� d���3���3�'>�8!�f�(�@ ��-��T��/��d�(6p�@��M��b�R����a!���MAT����Ñ1��u	�7tMџ4D�$�R���c/J[��y��C��y"�7���#�m�%:���Ѱ&N"��'�a{�*�Ȉ��Q_r���/���hOq�p����!��pFAsa���
	�!��B=g=�p�C �Ct�)�٥N�!�$Ȳp��D�_08��a��cw!�DK�o��m�tEZ6S�L���>7�!�dΨB�<�+X
B���t!�D���"l�E.�'*��X�,
�{d!�� �y�tJ�J�8���(#E��@0��	k�O�a���u��Tk�>�B��O>��A��Eك�A
dr�8D�~�,�o0>WQ�"|R�'�呲AK�Bj�����N�r�'i����E /?�-:��@:�MP�'��i�jP!:d9������'7��� XB\���1R\��8�'[O���?�X����<4�``���"o��y�Cj�(8G�IF���d�$�&E�p���F�l�J�k�L<RA�O�����	f �X��:_�I(�@H!e41O 7�.�	���'?��&F��x�ycP�*E ��� �	F�����)^��%�EH-@f��C�I�S���Dl+_�\4��M6?��C�Nl�����ݪF�� DK�<�nI��'�K9~kr�C҇@;e!!�Ak�P�d(�S�'L�T5s3@�<u�����TRN1´�)��LS1@��~�9���W�k�&l���,���<��I�.{bX��o2Y�X�a(P}�!�Lx�|���b�6QԦ�-L���s�yh<ٵ�.^H�\ZA�\��|��*M�<9�!�1���#c���'H(F`���>ɏy��.(�
��cCQ� T1Ak���vB�Ɍ_�J�QoS�Q;r ��-U�t�V�I֦�Exr�C]RZ$�A�>�z��2��:���y�*�#(P�rT�=;LX +W��	?�V8�ȓJ�։Bʌs<��r ���T��	d��hO���c��z���^�Y�bބ|bB�ɍK�RԀ�s�)�G�1	�B�ɷI��x[�.��2����V%�2�C�I
4�؈�r#��y&�8z�ӻ?�0˓�0?�2F���T�W,�}��daѩ�iX��mZo}�灊G�ޅ�Sl]
e`�dr����yR͚>y�����(`'6��!�µ�HO��ڌ�ɉ�3v:\Rb,
�B?"�3���N��B�I4ZH\�G��<f
�ࢎƌ`6�DK�������G�9!�epu�	
R���@���y"��#!�DM�"g[!谇����y�
�s�⠣��Ⱥ 9v�F��>4���=E���> (� `��.&u[�Ν�G�ą�7aV�	ENU��$|rB*S>"'����Ȱ<)�'��D�� d�P (��s���;���,%�d;�O����E�r�r �!�*R�XC��'A�OZ��+$�
����Y�n9N��B"O&a�'d��浻u���Z@LA@d�g�Iay���'P�0 ���;,J��t��$��80�'a��oϏ��*1�S��J���'l����#q]��͌�R��¶�_u��B䉾q�ĵa��Q�̌ɥ\%d,���v�xI�D7.u<����*Md�l�#������J~&8�7D�<T��7)R�~ԱO��l��H?��-;��+e�(I5@mㄊʠG��'�|"ŉ�/��`!�Kϵ�ޙR������$>ړ�~⅝�����QERs<v�߶�O<�>1ݴ�M�C�I���-�6��x�rTB�bRZ�������:o�ܑ��˄�h'��Y'H
�wyfC㉙��Y-��Dbb��l��B��hC|<��D�w����
�S}�b�D{J|j&.X���C��?�V�0���V��hO�O��m��'�8,��%�$�BD{�'pF� �ԏwʦ���)ۓ٬��'�j<�a)��_��$Yē�Gv�R�'�"�
5kX�Jw�`9H\PAi���y���Uz��yS*ʄl?m2v�(�y�)(!��a��̇cI>�f�8۸'�ў��� b��j��*��
�x�X��úi��	I�)��q+�O(=�܉�R7>	 ����8�	y�$�/�(O�N�;�p��v�E�`^@8"!�o��O���$��i,r�E�ͺG֐���: ��i=��'���?�����D��\V��Z2���,RQ�%d�!.B�&
O����],$��v���5�U�D\�hm�h8���F+P�&�x��V���{� ��;��I���Ө����dFI���sEm�۪˓�hOQ>���NL�3f�A�N\�Z6�ܛ�,�v�2����!*x
��6�vx�G�aZ!�D�16�ΖR�&�nX-�X��'�ц�ɑӖy0��*�
l���9<HB�ɓ4���A#�
 s��E�N�.B�*��@8P�H�E���k�2�
B�I'[�"��]�B�e*BB�wP"B�I3L���!#x��� 0l\�VC�,mfEi!,�2��H@���K�HC�	g�@!oV�>����&�W�oOC�87���oN�b����"DT6L�C�K�b�@�	a�@<iA�R�TC�� Lt���&��&J��-Թ�C�	pVH�G��$T�0� �� OS�B�I�|�����́)7�HTȡB�}�C�I�>��(���<8���JF�Iz�"Ob��5(-�<4zqm��
�,��"O�ce�w�T�c'���kf���B"O�'�Y�G��s��ǺNTs�"O� ��Ǉ�
� pv/\�
 �s"Oz�j� حr~޴����H�����"On�eh�B�&��sf�&Gv*�CR"O����mݞ	S''��(}j��E"OP}{����>��RLY�Po�$#"O�i2���!�q��V�:;XlP�"O"�(uA8����f��	��_G�pF{ʟ(�8ce	3^�Bm���G�>:B)�`"OY@��T!A��i��6}��9!%"OА�FbrD�&O�q��٠��'o��`�d��G�p{��D'H�.� F��!�dU$��ۖҬcy0��gD�[��	{?	b�铭2��H�&Js�0Ҳ��]ÂC�I8<�^\Q�`�w"t�1�+M�&���<�˓MR���P�G +O���p�10!*��?�TQ8�*Y�lA��"�0���ȓV> Q 
-"\�z�d�-�5��&�
�hV��W�F=����l�܅�_a��H6���=�ȑ�dA=
 �'�ў�|�Q�WS�}ҳjP_����¥�m�<	ҁY)X�!�׫�6|�8��%�R�<�܄&���`�����$1���Ye�<�g�Jն]�`i�"���k�(�a�<qU�U��n�s5�ӡ8��-�"A�X�<Q�S�Hc�i�'�R�!��	l�<��n-}�J�b�ƍ���ę��]�<I%�X�5z�AÏ0 i�y"-\�<A�R��hQ�7�#RHf�X�<��#�3h��8��ٶ=E~I�C-D�8����-s�q[Ǖ3A�B�2��)D�ةdOW����w��!�85�"�<D��p��R�4�MF�.*V�:D��9�Q�h'"|��&8�(�`�6D�D#2����dtj"��>M�yB�9D�<RWc2,�2D���\1i����6D�����N1Z��7�کp��8C7D��R�ą>R&�rv+X�?��ce�4D�� T9���X�&��a%ӠGe�"O�{�ǶHxN�k���w>>D"O*�1Tm
�\(�1M??%:��4"O���❘{���@�Ⱦ:��c"Oh�ӢmH�>z�iS��JC"Oz=��:SY���HT%*� Y��"Ox#��
`�ib�K��Z��W"O*B�o�	�@I�Γ��a��"O(9�R&��h5k�Nk��sr"O4�S����`���QΎ�rXR0"O^�(��ֱ{.�pp�-7�N��V"O�q�g�؃F�(XC��@��ey�"O��#�ʊ?���G�I�8i�E�6"O |�S�܂_K��4N�4Z�X�"O��hF oRj .R�C�Mh�"O���EF^"��Pmދ63�B4"O����AN�aS�<*��%2"OL��BV���y��H���1�"O:Iy1�ͽ/̖u	�,�}�P��"Oz�ae�ȄtɄ�1��V���27"O�|��k��@$©��/��W'�+�"O�Ò�N���",ˢT����"O
<)Sn��&:�#���(�b�,ψO Q��K&)$�[F��|��E3OX�y�f�2m3�\
����ޤ8"O�L�� �2F,j�:���!�m�"O&�����z*�p'��6>�-)"Ot�J�i�<_����B̾]ԴT�"O�����E�6!0-H0!��.5i�"O����5]!(���J]q��3�"ON�`���	G/Fd�5N�;L� !�"O�l��D�)b����kI�	!�ؖ"O�<���f$ �	��� x�u�r"Oe�G���5r)�&qBv��"O��s�(�<5�k�U�zڶ,��"O֥jF+C8]
��t�8T��ሱ"O�����B1E�z��1ʊI�V�@"O��#N�+_v�����e�lB�"O�UDjI<�IC�,�#'��$"Oe$(ЂWJ��D�F6;�X��t"O�	k��	G�N5��?Kᒨ*�"O�d�Ac�7Wp3�(�#��� �"O��Ї�Inꁐ2l��S��8�S"O"��т�9c���F�P�U����"O�B�ŭBS��w��8X\��3�'YX��g; U"��m�K�P����ڌB_��"O�Q�E	jwB��@��~㨰5�	�Ң��T!�: �t��@��?=uI�HX7"O^�p��Q�&E��N�?A����տ �#E��5��������썢 7k+ ('����Z�S��B�I�JP>U�7�֔9�(m9VLͫJA��������)J�flV]�剸 4�Ëa��Y��CI7&������&׀+�n����dZ�%�����¼N�t���/$�s�Bŧ+�ļ��:����$@?�L�-��-�ʨ��4��N�����NA��2�:�y%CV����	�,4o�8YB�$P6�X��		�h�z�Ư<E���}fJ��%�ҫ=Ӹ}ieN� g8e�ȓm��R'��<(v�U�`gޡU]v��(��a���[>���
�r���X �ԘQ��$Cc���U/J���ɵ3�Z��n�k&��#�@B32J<ኳ�E� �ZE@%"O}H<�`�ʕr�6�; �'j� -�q�l�'�`a�E
�A����ϒ�V���bֵJ��4P��C�<Q��XTZ(yU΁�Uk���G ����e��V�L�	�}��C��[@�O E��0X��<2�<���ED�!��B9�j�Z7'W'E��]p�'.,�&���֭wqp�'Yd#}֧� *�u�;4�:�@�� �ls"O�L)�9�-Z�J�z[B��j��3���A��F��̄�i��2�.�.R"�S��|K��D�.r����0�	2
��IK�{���oڎY���􇆎'��l{�������$X�=1~(	��[��� f�B�I�-çA�\��Ff��$P��\ÎT.g {gB�j�O袤�E@�<�����(�;�1�-Or@.J~����G1G�a��̚%VK�<[���*����`
EĴeEO1v��ʓ-�|�'�
��.-&�`)�� BOl>���h����(���f;��$�bH0�"#[E�@5��Q
�B	���->��T��s8�l"!d�v�x�·ڰ<�v83!���g��}
7	+y�G}b�2h��)�Y�r��,e1����	��,S��	(�E��8�s�$f������S%�Ksn�����1���D�5&ML�R��֯^�Oa��0��ú�8s`�P�4��q�2��"�:����1��+#J\��h���I�*�jE t�JBC2(�I�eY���@S�p�O� E��O��N�4y�z�Q�f1$H��V���y�Y�G�wh^	"�	�do��x�'ٞ�CTN�6"�C��
"��i���D�a3RN���(O�2#LY�!��q��M�;G~\!pϞa�����I�u^�G����SVYTm:�����D�[@Z0�=Ib��/%'��0�ȣk_�up%E�$��Z�19�i׆(s A�)s��ȓ8��E��i�,�p�X�",8���ٓ+Z����bkW�*�Ȓ����|��)-�r�'���w9��x� T$ʆ��Q�R��{�,X�XK�;�9O��+qc.N�١���N=� �֭=0 �"D�pq��30��p�kY8[�Ā�"#�NY	�>A�!ӗE��ذ�e� :s��� U1Tľ82����ƃ��0���?
�����/4�4%�?:d-q5G̓4�9�bעU����S�V�<Y��Q�V jJ���>8 b%y͟T�λW��%�d�³0���A���xN�,��'1b�)_�-���#PkM�jv��B�#F���b������ͺk�hѥz}�L
��@m��nή��Sc\�;T�%A`.MuAd��Ċ1'ԙ� �ȍ�?YV
߉+�l42$΂��f�q�e�����+F!G�<(#�Ζ�����D��K��M�G��9Q�>D�e�^�2��O|M�w'�%;x ���L	�`�֧~w�L�S'R�B V5�S%
�<E)e�X![�Ȁ	4"5����K�� ��7y0a�F�J9�x��4�����҆��/ٞiA�b�:�d�i6d�}�djޥ�C��u�v(���	~��y�+D�4	v�Ҕ#n}�3%���x3TbHdL:ii�`��8^��ka��1A �֝KV���	��i��'?1 �m ��d�@T�,�b��T�����,R�I�ɔi���+���$*�ːEG�Y�� M?|��mX��L!�Ex4h
��G|� �Vf ,SP���Oچ�qу��OxxST����y��R�]��%�#b�4C[���U;g�`� ;������U-V�c!FO�\s���䜌U��۳h�as<���@\d�'r:�¥@ݖa��0� �9���)F'C/\�A�O:�<�+J�����͐�|��9��'I�$�4=���OC�~~��0��#Dhy��O�[�8ԩ�ۑM��>��C��Ƽ�6�Ѵm�$�i�D0w��԰dn}h<��ne���p�+�^g�QzHp���	Ϙr�Z]��ڤe�|a玝c�#=��̄8붐�0�P���Xp!�Nx���@�Q/ ��| ����@�s�(�.�2��(_@�<("!�U��܊�n�22a}�+Ãd1�h� ��6��
����3�af��h�*(��̗�vd�#��c��]����`�6"���4��4>7���G|x�5FA 0��H�,&"(vh�ɕF�BG��I�+*"<S���T��]>;&���IEY��1�L�y`C�I�\�Έ�G��FTn��Ã�^��u�U��y��X4><:d��*��]��7鉨''�E� a�>h*���o�':����$B��^D{S��%Mq�3Ť�<m4�͓g*�Q�l���ܩ�f�d�Uːhx�xh�Bײ6�(���ߗb��+4/}bEU�,���(О�R�J�F^UT��r̜q���ӿzPB�z0Ϟ�hK^*D�yb'�<�4U���X?V�����a�A~�i�l_���s%
��j�mK��T�4ٴ�Ʉ=ȱ8qD4qM�IZ�+�B����Jf��s�J�HV+؄��"�@�ckA'��5�d��ҍ�-�*��$j�U�g�X�Np����My���ޠ`�"��#��#6T�u�3��z�`�feI\|�\K��O4��9�Ȁ�B�I�0?!b�GhZr�a��>U�$�`-DP��_�~(�T)�!�!F��0s��/8���B
�����@-&�pc�ĸ�B��Ń �q !�Y�2|5�'�K2�ɱ�B�1�]0pC�x���W��~'�xh��	��Z2�A�'Hh���J�z����E8P�`y	�'%0q7#ԓc)dqC`Ö�k�4�э�q3F)	��61x���O�� �@G�Rħ� X���])�@\a��T5_��c�'���艫o��=�g��,l�֣P)7м!�ƈ�+I�)k�%̈́i7�BC�;�O	�d�&��x�V����f�|�L֐��݃��P�I�(@:B�J6�l��?����͖��| �&U�"���Zv%}R�ͪG�;��|���ݔG�p�02@��TFP��
�q��&	����D�*�� ���INb?���)P��%�Ő]A�|ѳ���#���'������]���Ϙ'bB�z�י5�����״&�\�2FD-Td�9SO�_rUC��,2bF�<)�ĬW��iz&���H��[ ���c��Z'd�4ɉ��#�]Pɜ�4��eRF	�c�\�V�É�X�B��")�����*]�Z� `F�T����,m
l�
��N�1�i��a�%ڸ'�0��@#�,U�baC@�X�O�4P
�%�XH:1˗(���.O�p[�i�/Y�LH�Ç:�|��t��7���G��hu�bB�)H���xK>B�>� C<+����c΁v��Q��M�
:̗'�Q��-K�n.�ϸ'CD,kt���� ��7DK;�Z���F�q��* \O�)� }�^ԊSF�3�� p�
C�=�
=��o�/;`�O9��O$��?	���T�|��"M�1t68#��.��6\q�e#
68��A�ȟ����ŵ;��lA��/�zCq"O�,򒪝nkJ�Т�Z#�x�_��9�Ki�"��6��~>1z�MY<o+$u	i���q��F<D�̐��=ݨ0�G�5�Z,@���HiX�pR��y�g̓m0�Y�Kҕ!UT4���-c`�8��(�y��=e����� �d��d�L��Z�[��p��͙G��	/�9��G�q��Y��DM `��B�o�h�C��_��<�ȓ|U�m8�%��6�V�T�-+؁�ȓ.g�	H��W�8���J0H�+��5�ȓ{�� �t�
�&p��,�_�2܅��N�E��y	�,9e��0�e͈@�d���}7�y+���X�ȁNU	҈d�<����S�8�|#kS+;&��6K,�!��ߚ =�$���C,00���QF��8��Ɋ!Q�=r���L�^`��gݮC��C�ɓiV�i���M8�t̒`�5kD�9������ݦdf�xI�)�Hl��	r����;4����<�E/L,W)|���$[p9�W�F)��A�h_]�r��<I���)�z��W$֊mXK�ȓ�S�!�DY�
��y��o�rld�CN��p��I�Df䴻ԇ�8S�%K�dʞL\>C�:$�t`)7᜙4lE2�� nLC�%n1�	�逎O��t{��ǿR;,C�	?5(�s���B�'�|��33D��
�`^����!��|�1D�3D�P�$ Da�9�4��>k��DC5E#D��nm��0�����9�Ĩ3<D�l�����WpP�aT'�&aB8D� �FG3S ����Q�t�JA@4D�L���N������eU�t�tIq 3D��1c�@�r)N�Paeж2�^���=D�,#�џϪ�Yw�S�|�P�jC�>D��q��!Q�<�QQ ��ExQx�A+D�@k��J�.ٰ�BȠH��Z�(D��Y7�f� �p�6�y�h%D�xP�aåS�vaҕdρ2�D1�"D��K�oǔzx||�6)oV���2b'D� �4%:Mm�X�4q(��2K"D�(��aR�_"U�)W�]%4�g�"D�(�w���0(��yw$�%5Ɣ���%D��0��]�$�cpOۗ4��l��<D�����:�� ���S�ʃ�'D� �$lU�h5�8��I��̂U�+D��3�'����0�({�����g)D��!��-!l�0��Z?���;D�(�1��0>��[6M�y���Ӓ�"D�� n�z��_. ��a)T;K�� �"O���� ?���krƇ��<�Q"O���,�7��r� @�DH(V"O�E	����p>܊�oL�l��Q+�"O�,8����'��
�!p�|��"O i� �w�m��.K*K��)�"O�Du�Еv�-jǈ��k�V���"OB|QbX"Gxh�#gL8�x}k�"O�t�T�/~�r4¶f�/Je�� "O�A���Lz8����s�֬��"O ��g�ÐahL��ԍD?5��0�"O4aT_�E=���Ц��R1b�"O����(��0e��D��X��"O>�y���^�mC���Gü�B�"On��b���m��
�1-b5;�"O��i�m�MjX���\6��a"O�=��-\��q���p�NI�d"Onp����	;�,��r]6y�B��"Ot����'T<$�3�jO?�"p�p"Oz�k3�Z�2׾��4��'�ns�"O|��B���^)S�%m�9�"O��B��ZZ�)��U�(h���"O��*�)��u0T�uXN�P"O`��5H�=��u3"�?NJ��ʓ"O�9���
P�&4Y��E�;�Lh5"O�Z4&��oĸ=2_��E+͵R�!���� ճ���(���1��	@^!��
j��� �$\�H�6Y3Q�ܙ5!�$D$Vj�p��� G�*�3���;:!�$D�H*2
�K�Ys��
!�C�!H���sN�J��
V!���)]���a޳6��Ag�X�m�!�d�0=�!`���"�!�Ɣ'v�!�f�e�2!E�0�����K�h���ȓg�D��AF�Q��$�p�Z�X���yI.��!`´E1G)(@�l��2u�qj1��vU���Ub�(^ ����eg�x���D$��H *~E��2�N9ӌ �(@�0�V;o�M��?��[����$�jU��NF4��ȓq����f��Ļ�"��pB��ȓQ3^=3#�"Ymz�3��j┆ȓxL�-2������3�d��za�ȓC��q���HY�D�V�. `�ȓ,TPATJ�M��|c��Qv 0�ȓ3C(}��Cý\�VsG�Չ�"��ȓϮH�P�@�9UD� .ɆG; �ȓun����`�+5�H��%�%m�v���%l�rI�FΏ]��$��4CN�1�$�M��l����ѷ�ږOc
q8�B
W�hDzR�  ���s0-�g��;�-�T!��S���rgؼ�`�ȓj5P䠷�Ǭj�$�+ ��e-"�FCy�pВƌ���)�矼3���3�5qR���G�	��*D�����@�1o����F�9=j�"f����Yc�/-<~�1�qX��h�&.L5B��AN�T"��U.2�OrD�$nV�N6�����T����m�"cl`@$*Sh�:B≑vظ����*!W�0�-P?IS�<�d��pנٓ7
�+��O}���P��<�ֈ�"$,hZ,��'!�e��T�-��@�a(I\`@��B��Pe�"O�����S��?��
��m�0�Q��U�z%���~�<a1b�WD4��� 2�P�'�x?�bbY�K�����9��<���ީB:Vٚ��\	<� )���C8�@��Ȗ�_	��'ʓ����������ġX!�8��a>�9���R�VmxY1� </}��=��؎oK6��4�5�3� 
�Lي	�2���E#@����"O��J2fx4Ԁ���0b�m27�'��(s��9[�Q&rq�����Y��ZE��^v0���L�*�x%�ȓyHqS�͘-��S�͌�w9��$P�'҄�J�b��Y�,3���;��U�Q�A��1k��+D���h鬍��m^$F�d�B�� *���.�J���H
����, �2U����J�d?�TH��F�#��:s1��*E���a̵1�#`���!�	��(m�)<&��j��'�H� �`�j7J�O\��Ō�+Qd�H°l��el�)���3��$3!�ܮe�Z#}��0,�Ry#�㚪� 0�2o�Ny��Џh��;� ��`:a�TJ�	�4Qp ��Mt�1s� S�x�T�˒�G,�M0�|�'�
\*R�Z 91aKǣ/�h����d�]Pl�8�=���\�E��ҲJ��-�M�􉄛R��=s$��#+���"�Pd8� ����wI���F̡_�ΰ[r7-WT0WdA�~h�F}�h��!�Y��E��sG�vW~�Z���-,a�P�&�� ��O�5Rq�:��az.8zT�t�X�XO-���r��fܓRtrM���3����)P�aBb��ӥ�0-r���OZ1��	d�<_P��G_3L�)9s�S�<�� |�vu��g�DՄ &��N���7����7�H��	8e����I�������^F~�c�I �R~Ft���+��u�Ťv�e�������?ξ��-ª����?�d�ü�dEy��kX����V�k�n�YԄ̓�j`���:8�ni G�FJ� ��FV��X4M�9��↋{���ر`1�I=CHj���mt<� ح2T�L?a�!�� �(ms���zt�c�.D�Dr������<$� 舑��'k4�p�.B|�S�I ̤�S�����T?��'��b3 �O/��2%Lӳ~e:�IߓS�<)�&S�y�c�|:X�a!�܎VM�0�l^�v?��M��P��(lOI5�� Q��[g��,�Xr�����X@�U��y2�]$f���3�a	�@��߀h��B�lS�}+�<B�	'!�$��@'����5- 1�^ЫG��w��扙Y�(P3o��{��|�?�pm�d'�uӔ@���ٱ�"OdA���ߖ�(���Я|Y:̓���m��YiqH��Z��<��+|QV�0�Yֶ�#qh�[�P�h��a{B�����c������d��h�6�ۇ��l�m�f�xӘ$rE-�'z��8�	ߓ^��(�~dt;H��0��>AJ$
�bEb�$�>�Vj2S0i��O��a8�!A�{����! �/�!��W�9���!`2�^�Ǡ�%�r���Ɂ���'H�#}�'�F�Ca��i*�H�P�u���Bn�<��˘B�A8 �S;1���eGV��}	H�� �iz7�'�DLB������A�K@�/j0u2ߓT�@��ӧ�yRm�j# 8Y1cQ0��ŢH�נq�B 1�I %��O�kPM���O,	1��_��B�:V�X츑�I�5�Pr�O�,M;T�P���E�O�y��_4Lp�l��NXj!��#�J�e�$�Ol����+�� �c˜��d�(Ğ|r�ܩ�j����=�����hN<�J0�O�gG��b�i�m����%�dՇȓ,�HU�"��'pi`eJr�P(S��	�҈��G%tohmj�Q*T��9�R�i�(n���`�b�萅_�;�a���4z
B�Ɍ�>�@S=3$�9���8��@�J ����ß6Fr� ��8�*<�T�ɼU��+H��`�PJ?DD���dX�K��\��=BK��c ��L��g+!��B���2Z�����OlunX�BB9�O�M�T/
��"�c��ya!���|���|m
��߇H�����*W3|�g��B�����v<���%�I0}��O
�yB*��/G&���O��(G�Q������$?4f̘�dII�vz��j8��98�j�̻k� Y�� ή!�:��s$�;wtB�Ɠk�
�!��KAb�<��3z��Mb0��M�9D���1���^�� ��d+�,����T�1	��J��W:�H���	#c*$SŊO�u8�X��ҿ\�Q�"��&��4(7D��oL��2��*'R�p2�'��p�ǵŉ�� d�"��K��C'C��Q8�'W/�=�qB�9s:P��?��C�*=��q)�I� `��k,D�(���X�PmA%	'm0*5� 0}*�IZ0u�a)��q��јT��J?��
�h2�K��/��p�*Yf(<� eLR|U�%C"�t͜���h�`VR �Q:`һA�������Td#>�E�y���RR`%��=Q�-�]8��sH>� dJ�d	�>svB�^�a�L3��:$�Z����%q
��J��N5-a~r�� ���K#S�1cPa� B��&8dҐ�bE�(�j��q䓓pn�P��&ͫ.�3� T-{�)֙S.�
��U�Dat"O.mpA��Ҳ��B
�V~��S�E|�ȁm�/�$I������O�&@��`��<)��ݐs�Zy�#Y��>�8�	�\(<���%Yxx� E�� ���b�(�O�(a��'ǉQ3�q3 �-���d��Zv">��c�8i��s�A�:LN Hv�VJX�ly�B�;v��P��`�8��!.k��t�j��]b�EGĔ5�2���0?����4��W�Y�f���B��y�	�g��ۂK�:	Mx����8sB�y[���y���?�,����dt��ƩL>���//�*����Y�)�ӹ< ��UaN�1��)��l�������\�,I���0(*��&)?ʧm��d�P7TUʱB�<7�U��҆g^	M�<����$�>b>c� �vzSz�0F��)̴��˄�l�N���%F�`�pL���[h�H 򤄢n�@P����U�������6d�&b��Uy�k*�]�vH1���c&,X��	�3Q ���\���K�����&�9�|�Xqw�͍r8x͟8��"¶r���!M}�z�q�>;��;��D�����I tDh��kW�I�H�IF��(��	/_�2�CE��O屮�ᓪ Hpp�C�EĨ�����"L����a����'��#}�'%2��b�wcZ���[2g�b!���S���䛆oÄ��u�;���P��Ȳ�:,˖=��.�7���Y�-Yԩ��/ANl���O�.�d�؋��R�!�+~���R��`��0rToܤme>���ׁ],�ړ�1��p�����&�5YZd�̟�8��O�j��1��ʋ[�T35"O�8pRN\�{���D)�,y�AX������$_��Q(�Ga>�P��'�V3���(*R1���3D���c��jHF�	���Rr@,��>��	���,ƘϘ'aBx��\%T��X&@/����' �e�i��ݣ�ah[谈ׁ� �����'��1��Ŏ�oI|p�����{���'k�݉eH͞9l�9��"�R�$�'�t�i�Ʌ�<V(�� o�d?j4�	�'�^D�w�Ү�L���(YZQ��'	@�V�N#(��jRjY�'�V�񣝞n�I�W�O���B�'�B�n��q��)� L29���'s�y��G�.N�jע�	5P��
�'�Q��l.asW#U(]a�}�	�'mƱ;�ׁ[�������p 	�'�8�-�(j>�4+$k
�r��  �'��ł_B�R��Å�2>�0�
�'�L�)%��b�c���+��)
�'�\t( mō8��[d	\�6B&���'6���H�o�Ԕɐ-�xJDh�'���`T�2,�����3{MJ��
�'
��+0CK!}��W/[2���@
�'�*@
�H��������ڼx�~�J
�'O��;�k_,O�
��`���J���'kH��G��^��,���9`�Q�'ւ�R"�
�]#���4�ԌC��	�'��A�	�1@�(�H���SKଁ�''vܱ�]� o�5���YA�ܵ��'y�M���q�6i�Ӥ��H��C�'#���� S�8��	��.	�v�3�'G�A`�Eo�Ż���s���
�'�&QZ4��P�9�f��i1�)�	�'��p�GZ�k [֮V�^ ��3	�'f&)`+�X��ٲ�i��9֤4r	�'Ѽ���F�X�&��u,�>"���	�'[̔��c�Μr�
�ݘd0D�t��͋T�L!�p�ʡ	.9V�<D�����R�+�Л)R� cWm��y�@�����12F�< �LP�JH&�y�iH!i�x��S�YV�^�cf��)�y��ԛM��%H�6IY��y�"޶-m��[��4EDJ!��'�0�y���-�>T`Fɔ,Bl��	��y
� �X�Є�529뷢��Q�옂"OT�qUɵa���F��+����"O!Y� Ð��ia��G�y���V"OB���$��4�`ꄯ_-�Xa�"O\�K@��V� ɓ4k�5�%�Ύ�y�&��J�laa˔l�2��T��;�yB���w!�3bU�y�%�9�y#8��q�E�j)�,7F��yR	�ݲ@.��؈lY�
���y���| ��9�P���y�iQ�g��Deɱ��Q��N��y2h�]�N�S�E'>��}����y��T,=B:��WAٴY8�rL_��yB@����dj�&\:\s��w��
�y"�ׁJ�|t��a�9/+�m0Ђ��y2cъ-�~ݹd>xL0�		�y��d^�պ�/jHCFU��yR&��+XаQ�v���y¨�(),� [s��1cfL�y�۩�yb�)�(��vM��\!�y"b
<�|q�K$JҤ჋���y2o��mc�ɫ�� �r�L���B�y�$Q�[����OD(�N@�`���y���
�lH�5� �^�vlЁ�y�\ E�,�sA�E+� �B���yB�hP!�&���B��i
�y�aQ�-�����k���Jܸ�X�y��ͽ�hy:w��O�y�.ߺ�y2�/=d�u{U�ҲGЬq�d�>�y��\�|#P9aQ�֤v�j�H��ȝ�y�`H2��١��Hc�|��6��O49�5<�%9���dO��4Ok�W65F�U�,��p��8�O��9b��>`�f��H��}Z`�;i�p�uÀ�EH��)�З璸��/?Q6,�O?������1��01
`42W��-rј3��OQ?�㴊���d
u(ڨ	����O��=E���[�����	2[� P;5钬�hO��(��J��Q4a�6	�1�>Pj�i(1O0�S�O��%�s%��Xu<���P�H�H(O`��P'�<A�<�'(]-��b��ٲ�ـ�ĜL�\��O,4=�'r0aק���D�Jݲm�cL$HHE��AS�8��y��)&`�lH�I�< ���MĐ [!򄑮U��A+d��s6jtSacG�>!��%,u*)B&�: �u�����!�D �*�p\B�I�Bh*��q���Qx!�$A	W���2 �#KZ<i2�}f!����L1��O�L6]���zQa|��|�`�Z�(I����H��fM#�M��'�qO��N��O���l�TXi�D��m�����z�����'KV�Ж8Oh�E�T��̑0'ު(c�X���R�\"<�缟@�B.��ĉ����J����
)"M�D�����P`�32�x�����@��d�'�4+K|��C=�	�4C2�A��-ސs)n�c��L#W[L;4#Y�N��	1��ƻvh�4z���O��s�`��j�O�2h�"�<G|��8'�@Y����.!��{ԧ)���:�1o��Az`�aTD����,S�"�I$���Ve�i>�Ӻw� ��' �0_}>h���[�y"ۋ|��Ol�����cG� ]�Ze!�#�[L���
>wڍ{��#�: �"a��Z��d�s���-F!#�"O���	\�*�fJ��O� �"OJ�1��Å`�4��n(9�)��"O�!�Ǝ�=�Ļ�k�>j�ۖ"O���H�}��)c�JB�]Rě�"OE1�� M��R�c�#BTs�"O�%ۑ���a�e�#��`
���"OV��I�/r��aҦ!$
鲥�u"O�!�1�q|�4��Ǥbz`e "O� �t�e�['$�Q���+z��y�T"O�e9t�	c�1�D?Pnu�`"O��"�[�O���8ҁJ�QN��[�"O�@�(���ze��=eYJ�rb"O$�b�{���  [
TE�%�V"O�Q1��=�R���N�9j':h27"O���!��#� ��S-؁Պ7"O�m0�C��x`X�0vA�G��Kq"O.8��ۙo�����O�
�V�i�"O��2A�A�\���Š�5!�n�J�"O�ɻ&ɧ�"mHG 0�0�z�"Oe[�T�!�ؔ��ᖮ ���"O6�Kޖ��0)�!�!�R
�"O\�Qs ��S3��)Q��j�z,�"OhT���߮BX��jg��!���Ss"O�\b��Q������t�+����y�O�j���A��w=P`ᄥ	��yB��9�IC B�mp����W��y��Ǉl/(�)��mV*P�
�y��A�r�˔��s˒����2�y҆J�Z�θ#c*֪�䢖��y"�
�p��)E`��h��s�M�y�-,^��R1f^�����yR��=��#�`ë����'�(�y�G��1���b�-�5�'���y��_�'��8B���4 �X)0G����y�$��O�L�"��*A����f��
�y���`�LXjd�#�&�ҵa߱�y"i� Sg�d ��v�<�0%X��yr�_�qb�	1�(��lF�������y�̎&�hB��O�O�V��VH�0�yb�UK�~e�Z�B|)0�Ͷ�y��C���!C��A�< �p �DY �y��d ta��+�*l�U"��yrd׶#K�b��*rD����yre
F�XSl�4)��ma����y�a�:�5 ��r�\�hT4�y�뛪8�h��сF�
�Lܩ�H��yB܈Mr T"XQ;�@��F��yr�Yo{�a�t�ٙKy2��
�ydZO�x�+wY)8f�������y�-�/W4l{��T�=ؠ��7�y��h����n P��HP��N��y"��0�����'�AL��3���y�m�r��2	�j��SC%1�yrFV=nk�ac-X�l(�tAb T	�y��I�EE�P��iO"�Z�̄�yb�ӹEd��$��9fT����_��yrQ-B�j��1 �^��b0�û�y����F��s+�	M���j��� �y"8�,�3�@fp��8�yr�H0U��az�i?4����Fc]��y�;wL@��Ά2�$U�wM��y�I_%Z[���aǡ"��w!�-�yŘ�Z�A�g���!�*X�6m��yBӶ{��T�Bb�$.3�ћ��8�yBE\b<20���N�y�P�U
Ë�yb�L~(l]9B�1kH�K��Q��y¤�D�����Ñ{$��Jd���y"jQ>6��S ��<+jm;��\"�y"eC.00�����D�:N���qZ�y���)���X��K�C�H<���;�y�L�J�8��O2C�H5�w�P�y"�G !�Н�e
ˌ
ִH*��א�y
� ��꒯�2*�b0��ĩ0Q���"O�4z�!��q�\XR-Ύ6��{�"O�d���E���A�A͗�	(<X: "OP�Y`'΄E�
"F�~����$"O�5��ơ��jڊd���"O����B�%<�s�I="�Q"OrM�PQ���0�)�<��"O��a
֩�~�EJ�s���"O�!�\(q�T��GBa�	؀"O�e������ȽQ��{�aI��Pc�<a7@Xp( P���l�h��i�s�<Q�a0�fk	�*ٸyk��Ol�<��!+TX�A���K6\]ST�h�<y��38hl�LZ�F�>�Xu�c�<)���3B`����� ��1�%�x�<q�jܞl�Z�7
��b�ↁ�o�<I��E
P�E�t/߲��%�eBt�<1��,K����t#�X��0��Cy�<y%KW�>��9s��
g�5���Fs�<	����c#�I�%pa��Z�<�MDl
K{i���L'>�B䉟� h@`a·PIz�YcLG�/2B��I�PP�amb���Q0F���B䉲$ʼP4��!<Fڀ���5*�C�I8�|����*+$�����0?4�C�I(�<m�!C݆87`�8��_�!��C�	9v�2�� ��z��Ł����AϘC�	�"�X�uU�K)�1Y�Ƌ+zC�	�(Z(Uq�����)��aC��B䉮OV\-`�MM�#�X�`A;y#B��N�TSa��l6�@$ *V��C�	8 F�ʆa7aP�\�%@:F�`B�I>.41�l�?!�h�h�@�q_DB�I�@=2= a�\�7���G�TdTC�I,rE<P�#s����g�&�DC�	�i�ʑx�d��r������C�	.�88��(�7{9v�2B��*)�C��0A��c�ps��0&��2ޔC�I����6��[orQ	�I85d�C�I�+Q*ps��� �(�@����VC�	�	�NyEE3dS�iǡQ�0�VC�	p) ����8J���O*Z/8C�%�>Y��H1����2,͟p�C�	�g��Ԫ�Â&D_Yc$˒c?B�e�*�Z��F�e	&y��a�B�	�.=�`[��1B(D�����#��B��8S��ShҝR���aq� "��C�	�fx����,��{��m�0jCϨC�9�"����V�*�����(�f[�C�	�@�l�(0d�'.���e��I�|C��x:<�0�]�r��� b�Z<}-PC�I`��a&IH>+��3SgY�edC�ɚ�`�2��1T����J�hAB�:nl��T�,VӒQI`�V42��C�	��t0$L$�6)0�T
3�>C�	�#L�b�֭\�*�ٰ��yXPC�I�|�4;��(���A�όZB�U�2"��'�j�"��+|��B�I�U� xz�i��f����/��B䉣	�$-�Dh^ m �Y���fB䉺Q�hxp���R�̍�3$�17 bB䉦2cRA� F�baz�"A�P#�LB��'Re�� E�`�8�B��-~�@B�� ~b�M��'E�v�Z�HFoκ<�B�)� ~�*��IvH��Y���kK4ĺ4"O,�!���@��h���Sa�%��"O�]���3zh�(jrIB�"W���"Oƽ!#�.�,x҈�'V&��hB"O. نEΩU.𻃇�H���"OX��UM�yݢ�JV-�HI^�5"O\ԁf!��Ln�0*�0�v�R�"O�h�"�h��֢�2*� ��"O
E� 萫l�P�h��U]��h�"O��W%��k{"ɹR╄\�.�0"O̸# �3W�,� L�P����"O��@"�!gԭ[�I`v�i�"O��0f)�><:S��W�pb"ಶ"O�`��"��*���	V	��&`j)3S"O&4sw.W�'��0c��[P�"O�Hi����1b"��#M�L�q"O��B��2lJ��/D1hq�s"O&]+�����-)�̄4��P�"O�!sp�N Cb('���M��}r�"O-����$Q����
ϓr����"O����(�jEp�K��q�"OބbB,]jE�ř�$�=7�d�	�"O��#釖n0�IRV.&��h[1"OJ�����+=�h��c#���
�	a"O�88��R��i23�Q8h��V"O��w�H�"Ȉ*��'�(XU"O�*2 ��#�:�9d(S�Y�Us�"Oؙ�vcZ�}�VQ�W��3.���$"Of|���K���P!�90���"Oe��S�8���q�o�4%���!��!L9�!�V�V�S�.I�0��r�!��R9�x]����2��P]+ "O��Q��N4����ek��v+�8�E"OD��%��>�~�8U�	�wpē�"O"��"ω@x� ���_�q��"O\!��)J�3#Ș�	�е@2"O��7�"��s�Ć�S#؅"O�T��m�|^�Q@�L*3����"OPm�Ɣ1y9\EB�,G$
v��"O�hKsJ�*a ���LI�d�80"O:)ZC��`�>�alY��X(�"O�D�e�IA)���aO�=�81�"O�1�M��p�I��ry"({�"O�bF�S�g�.Xۄ�K�����"O y����2��t���]5!�t��p"O��w�l���G��[�U��"O�}��	 �0B���舼JVN��"OQPBl�4}�ب"g�._���kg"O���vޓ��eyC��?���9�"O�t�$N�)�$� �d !��Ţa"O�ٲ��*f3~M�4�Йc���K�"O��y HɠE�t�	��V�\�8�"ON��9t�Ash� C��y2�"Ot���$�`R�[C&߻q~�	�"Ol��ȍ�g�Uyp'̭d��x��"O�@�b��	�Va��'�6}��T�W"OХ:PCR�(��� GC1N���;�"O�[a
$,E���V!a9R��1"O~�z��@�O�Y9U�Z-�h� #"O�	����nn	�҃�<Q��<2"OH�@ 
  ��   E    �  �  ++  �6  ^B  'N  7X  �`  Jm  !x  i~  ��  �  ^�  ��  �  (�  j�  ��  �  6�  z�  ��  �  H�  ��  9�  G�  ��  3�  ] �
   � @# y* �0 �6 9  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�ou�!Dy�'�:� Ή�B�\O�|�����<a��$�+q��@rsI�E�f�W�]�1O���$���R�W����FޜO��'*(#=�O��)1�h�Z��K�`)����:o�.�<�J����<4���y`���`KR5��O��Dzr��`S��o[X�JC �+�lԛ�#D���5�^;Ki�e:	�L�� 3 �6D��@C�>y��HRc)ȓD�* �$?Oz��L�r�:M�\�H�| ���� d.���'�.���Ǒ����r�Hp*QGz�~RQ$X�E L��]O	�fe�y�<Y'�J�oW��`2m�V$��s��Any��'**��%�T�ncL�@���h���'���!#kB�踬�@ˊ	�2�#�O��G{��4F�R��F�|�Sm]�y2��6u��	��݆i����y��K�eb�#�-�b���q�����Otepa����+TJ y  �0��rL�C�I�t�@m��'[2H�U�LQ�!>Bʓܑ��|Zjͪ<\���,B�~�!�a�B�<��F��@��4�S�{hh����u}BX���ڴ��'4��'o��e�f��;i�(1b�蛞09����Z��� ��x	�aqP&�3^i^�Gz�D(O�e(P���0�2m����
ba���"O�mkF��f�-[����gX~��"O�Q��gX=L�(��kL�*mA���[ԟ�?E���P��,A��ޛg9(\���C�̄ȓy���C&�6��[�M:_�,T�ȓJ����X�%;4�҄�B�kTL���	|�$�8v��Y��l:n�뀣�;RV!�$ ֒��O]�6ě� �HT��\E{��� �QZ'���Ԍ����<	���"O,,�p"T]q������^`"OL�:���\�Pq��@Y)u��x�&"O�m�S�O)t�~T�%IM)n�-J�"O@|�㢇s���ʡ'K8IO�ܸS�'b�O�l
&C��~"��ᐙ;�fY���	4$E������}��p�'l���L���<}Bd!##,h@���W^`򣉒�yRN�C�y� ��"P��)��
�y��	�c�e�хI�J�Y��y���QĨ�J��43�e�ъ�=��O��~�ѩ0�IBա���@�@�P�<0�C!��8Ӵ!�0r��ЀRD�q��D{2&�r�P�;��O�_^�Qv�@��y Y,a�Lh�ؠden\����yB�U�2�C�iX`X������x�iNx�(Q�ԪP�1�C`@�p5��>y�'�R}��j�Kn�0@��G��%KÓ�ē5�����~YI��������d;6�}��!PdsI�b��E�3�\.I�����hO�>�1	 �p����ʚ��N�x�a2D�Z%mA<���Ec�u���c ���E{���\�d<:��$�%qp�y� ��!�\~�R'J��JT�cԦ<!��Rdbm��FC�^A(���B�!�D� &��59���XO"���A�)8!�� �Z�� �Q�8� �O)!�$��V���ʡG�=,��cOE�	!�$U�"�Z�!�A� y(B��m�+�'a|��V��mX��	� ��Qa�R4�0?�-O��ST�,��88�8H�
��"OZJ3su��sU�V�t�g��0$�,2ٴ�M�۴�Of�U2e�ԑ+!ƅQ�)B���'R��PK�0wxfK�"��m�H��1�4�MS�y��D�ȟVD��k�dU @�e�F���O��~·�8~X"8�aÆ.VJ�ڥH@y"�'���c&��*`�!��	x+̪>)L��(��Y��i�J&�9���~m
GN:D��C���"t���ԩ�'p����e2�I�~�O��˂?2p�`"�_T���' $��`�8x
,�S,��jl�<޴��'꠨�㉁��(	�N�(��l�eWSdC��#e٬][�N�h~�h��U�B䉷A�l��e�zVLaei�n��⟜�鉰n��A�x2THU&^�X�B�&7,`T�w�l�J�y��ij�'�M)tΉ5r�a�7�M61Dp�'�(�I�X�91�ɑ7��),H>�[�'%bаf�� �.��vK�:��p��OƢ=E��&�:Kw
ϝ]�
 �3*D��yr�ΆZ�>�wO�Y�9�ee���'m�zbiW�8\P��B�W@\L��/�y��R�*��
�2zB�t���7��*�S�Oav���?$8��B Ts�@�'&������:������/:����y��'��XB�EiRm��K��]o��
�'6��*�,X�� P`B��T���'Ax�oM�| �ɶ�A�TA4���d.�n�;p��$ܼ�;�KDu��Qi�"Ox���S��ϟ,.�~ez��b8��C ��-w���Gt�<Y��8D���Q�5$[�x��h��W�)D�(����V:��j����T�lK�):D��i���>������[bt@��B7D�� �t)�ȍ�F�!/S�D3���"O��mʀ*bfu����4j.��(%D� �pI78�ޅ1��t�cm&D�ȳ��O�>�z5ʀJŘXSF� �d%��ȟ����_�)7(E�KM�b�S!�x�'D��pN�:㞁��f�$%�j5�
���d�L����FL�D� x��T�!�$ƦC�&qb��@�(:�V�� �!�Dߋ{����6<��E<�!�ĉ�^�z���eN� N`��7�"f򜔆�@y@�� .�&u��|iv΂�.�,|��ȟ��OH���� beHT�dO��*t�ҝI��	��.�~�'���l��� �D�#s���'��l��] 5����╀e�Bh��4�~��'�����$ {�̍a�_��(�K���4&��?���MBx��˖� sbi�d++D�d����84�e[W�J6.���%j��O���ħ��/�v�Y圻��K�*��hƜB�	]袍cV��;����5�Z	dc��$�x#�'�ayb�����Fc��
V���w U���x2�ޟ.�H�3�E�Z���� �3x7(6mh�
���E�8��5��ǎ%nؾD2V,
�T��O*4���	A�uW�I2��:f��P k�j�!�ǕV�����F4$����I�!R��	�HOQ>��m���J�{lA�;���,5!� T���1��i�ܠ�M�*P4���>)'*B;F0ѡ�$�p�ڈ'�F�<�LU�Z_�H%	e��c���x�<��ϋ�I$t��cO�Kw|Yc�J�O�'1�O䠖O�h�O��j���X����h�)+	�'���A��"�b���*^�T�"Q0�Of����>�Ģ�f�!E4����֠i!�3C]pQX�N W>�i��a
�QP�_�l&��g�3�Ha�O���%:��тact�ȓ*$�(+t@2*K>�9�dܨa���ȓ5ю��@�4	�2�I��	�=�(i��c�����"���&���f�$�BI��%s����*Q�x�K���"5�^Q��:��Eɂ��0zGv�TK %�<��#f�i���
��TeM�kθ�ȓv� k�e�EB�䢔՘C�jy��)V����H�pE<-@�J�B�e��I�v� ƣ�
�=�b�8�Ʉȓ/�<ٙUn�
���u�K�XO�ȓd�S�+�{�	�c�%z��p�����e��Y��9&
�t]�I��P�� 1�(Y��Q���A?� �ȓ-��1Cdk��Z^�5�7�2u��Q�`=��NX$!#�$�&mC��Їȓ["4<����zO���&���M��V��U+S�0/bU@҃<7��p�ȓZG�ي&�^?�|��6>g���z<l	�V��$�Z �88Zh�ȓOS��r,ہf�ԣ1.�2fW�Ȇȓ.��-)��C�c�$8R�iäs"`}�ȓf�&<�b�
.^���c��%Jm���ȓ5�ڸ	g���K�����ʉ"6�P��ȓ5���GF�e��}����&Qv`L��:5�h+A��:��s���W{����qr0�Q@%yp-�P��o�&��ȓk�y#Re��.�ܬ`bG�5}�����}��)#ӡ� )E@�0��I�Go����\V�0Ň�e�Nܰ7dF�kԵ��%�܉����2�A䨂-&� ���S�? �Hg'��Jd ���3�=�G"O�a�#��//h��Rl�Y(܀�"ONbC�$�U�jN�J�kw"O����KP
M�`)$�Y;�"O�Qq�ʜ}P���g�T�ju�6�'�2�'Gr�'m"�'�r�'��'�048�̂#g�h�85
W�0>�d���'�"�'���'���'%��'��'r��g�<J���u��7�'>r�''��'���'���'�B�'�1eBϲ	;Z�jFk��(uڃ�'.R�'�R�'*��'��'�B�'a�a�T�I8*hⱺ&��4=�p�1�'�R�'$2�'�R�'}�'8r�'��Źw�P�mx"��Y�Lˢ�'��'w"�'/R�'ER�'�b�'���G�	S �]���+n�� #�'S��'>��'���'���'�R�'bP����F�n�fc7(�i���'l��'R��'���'2�'�"�'@���f��A�z��1� ���`�'_b�'�r�'�b�'���'���'"r�:�eć5����"xEC��'V�'R�'jB�'�R�'2�'���$e9
��	X���?.;r�Y&�'m��'���'���'���'1��'cB��.�t��1qs�ԧ%?����'�Z���':��'���'�R�'u��I�,t�+���b����ETjt�'s��'X2�'�'>�6��Oj�DX
)��X�B�?*"ts��
V��'��]�b>�b�Vk��=1�i�7�ڠ6 X�N��[�6p�Olmm�{��|Γ�?���Ϯ����@M�+v�̙�iĬ�?���<|�TX�4��Dc>=X�'���-[��`�F��%C�4PB�DL�N��b�T�	Xy��Sdp��� ��D��-�U��?o���4.��������y�O*
�"X�P��JǮcR杻t ��'��>�|䦅�Mc�'�La ˇ�&.$8ԧB6��	�'��d�ß`c�i>��	�٘$�1`�^m��s�»{#��	ByB�|�#a���{B�^Yj�{�J58R+��d����?y�Y�T����͓���7:}�����I>R�Җ�S0?���П��!��`�b>���'~����	�ƪزVJ�4�@���J�'��ޟ"~��L�:�Ć�%6�0I�hך�\�Γ+��ǆB�$P�Y�?�'*���p#n�� 7�Eɠ�m�.��?	��?Y1� ��M��O ��=��CC�G��0���!5x	)��H�6�Oz��|����?I���?q�u[�|�Tg@�?���B"�
xª �/O��lڶ!P�����h��]�s�@b�CÉK� ��?��rc�����֦��ٴYm�����O���� ��Ѐ��'P��@��]4?x��kV�ʅO�%���u���ڼf#��SV������X��a���<R�%`f)Ѷ,�a|r/g�rm���Ot0h��A�fJ0i��Ď�W��%�1i�OP%m�f������M[��i96M%bRX�0�ŽKbl��G��pИ��fpӌ��ß��g�K+�4a�Yy�OfW���Uh�"�#4�!3 ���y��'�Tᰶ�*J�J�sV��_��4��X���	$�M[te[G��!n�(�O6�Ȍ�zg�m:���^�z|*3&#���Oz�4�(\@�giӶ�p��$�
��C��}=H=ڳ�/���j�Ky��d�E�t4����z�p 'I?� �ٴĺ��)Ob���|r�$�
R�C�jZ�$>T5J�t~2*�>��?I>ͧ�?I��nd]Z���2;�� ��0P�L�@KZ;�Ms�S���S�Z���.�d��tʸ��D�p=6�Z�bn�C�'&�'��T*��Q��y�T�1ݴ}o
i	��T��L���]�IDQ�f�?��Z	���'��i>�	�O�ɷ(;=H"�_h�ٹ�o�"6l���O�%�""o���	��0z�@�:<:�i�<Au���"蠃���$�MSa���<�)O����O����O����O��'oz:��S�C;>�`��AL%d�@x��i��݂��ݣ3yB�'��dK[8	�b�'�6=�6����� D����0�L�S՘�;�`�O^��(�4�:���Oz�'�o��ɋb�x��"�3��0�T��9*�*扡_o�X1��O\�����<y�����d;�dh�*�> �� ��?���?Yu��d�¦���?�Iʟ���5$��ɳam�c"t��@Z�I�p��O,�D�O��OY�
G)6J�H�p�R��XD��<Y�>~����L��M��O����~��'���8��\ U5����W�8dne8�'��r�,_�SϮ1��m�C*Z�U�'��7�ߵU���d�O��n��Ӽ+�L��x����˕(a��
�C��<i��i��6��ئy�pI��A͓�?�2�J�_8��	L��0��ֳ7ԍ�6� "|e���J>�.O��D�Ol���OB��Or�8�˟bv�H�3H�)�����<�#�iL��0�Zk`R�'J���O'�'� �s�Q:eo��J�DL�}��1y�>y�������'��
M=��	�o��T�`��g�*��N"��	.<�ٺ��'D��'�Ȗ'�̈(�C�5��H2@O$`����
�J���.�b$�/aцPvkH�1�m�����yb�b�f�t�O����O��$N���@�g'0p��+��k:
y�Oy������4ruIG�>��i�<a��ο� ��`�M�|V e�1�H[���G5O���$��{�$��b��)���C)�U>Hʓ�?)�iI��ɟ�	nZx�I $<�x%��;�VQ#���2��$�P�IƟ��ɘSX0m��<Y� H���Wj�-�|IB<]�,�9c 'v�^�	@�Izy�Ă**y�e�^�p�j�
C/h5��h�4f�����?����ii��ȇ쓙�6=z��V��	���Y�m��4e.���4�O�R���獙b����A�
 Ln	(���ވ�塘\��	�?�bS�'op�'����eF�/Y�Lh������eE7�pP�4`�tA��Y4L�{�f��9a��� ŗ���Ϧ��?�V���	�e!Fx'F�q��#F �};X%�Iȟ�V��ئ��?)�F�@�2�Gy�C=��*�	։7��P��eF�y2]���	ߟT�I������ĕO�@��cș�l�&,+�'����4��	r�<۶��O����OZ�I��5~��wZ�����D	�e�1�Y�]H�j��'�O�)�O,��)��V�d͙64�X ��1��\" ��A�$���t(1��"�O|ʓ���W.,{,����O��Q�f!�Gaxr�p�ИK�h�<���$d�(�[<b�h�D����X��Ȼ>)��?�L>aFE~��3W���Bo�o.r�I��p�	Y��o��d��j�'��+M=C5r] C��"��6*�(0!��d] �GW��p��J+x�8��yL���%�r�'@7->�iލ� FA�r�-t�޼x��O�n��M���iJ(�R��iG���Od���&�*#T�\#��Y�KK�^���	�2v:-`v� M�j̀��[8�@ˣ&�lCV��E.�rU$�QD��&^J͠�F�Pj�!D��-Fl�E
�K=���'x�☱��ƳQ�h0XB�
do���Ʈ�O��� �_� 7�ɗt�T��wd�.1���2��6D��T��/{W4���b��#�$�4NK{�@�6���س��<P���m��氁�`��<t�0{���I�|��� rc.�� &	�] ��:�e�2�V�@ve��\�;D��	q��A��-'�l��/�R0H��Ƹ	�� /)�2DM�;G��5Cܴ�?i���?�����	�@��EQA*H��4�7��_	7Ϳ<Yf�^}���O�m��K�����"�8p��شT�h�V�i���'���O,O�����K�8���$8���{6�D&޶l�yU"<E���'/ڈpk
	O�����*f$%�s�|�Z�d�O���h>�'�8�	����1��]�$]�k]�a�c��8����>ѐ� `��?i��?�w�%�4�p��$� X�$�҅>%���'E6d�H2�d�O��$4���zD�0N�ry\(��ր|[L�(�P���g+�I͟d�I����'�~��/Y�@�-�4��#?�Y�E@�T2�Ov���O$�Otʓ�敻�nQǚ�pEZ's��̂*��I�1O����OZ�$�<� ͪT��IƜ� ��[Ĉ�J#(��O���QN<����䓸�>Wl�	�T�N�b���X��X��� ���?Y���?!-O� Ȳ��{⓸O���AH�\Qh��&�Ҥzg^�ܴ�?!���$�<!��N��OJ)j��֬)���3�@8`�HĈ��i���'~剔< �QI|��j�b��B��� E�L��& �@��'��	�,�^"<�O�r��7@�<GN�pY�M�%#��kش��\�!�=��'�?���"J�	 �x�q� �A
Qg�G,g��7m�<��|���OJm�%�+y���ɰ��� �6E0�4����io2�'��O��c���GC�z�8�W�ۙ5מ����M����W����K�Y>^m���u`�H��(�=~f$m�����П�)���>���?)���~b���$�h�A4���"��_���'�d�S�y"�'���'���P�ōI �,�&톖T�Fhpac�L��L�4�$���	۟�$��X�J����Į�Q�,P�SJ�2J�%P�<���?���?��O� xi�k� "����%.��I����O��d�O^�O��D�O�pHFE�1K$�Qt�ш��#��Q�a<:�G����I�����ğ<�ɱXl5�',4�!@�9u���s��R̤l�gyr�'��'�b�'��y ��ڴ�MK�F�&��y��!�.���L|}��'�'g��'��-�0�'"�'	6#��1m|�{���&7R�9��O{�@��-��OB��D&�T:tl�+��!Z0ɛ�l��y�fm�,���O$���O�xШ�O����O���럮��*�c�����9rl~��f �{�۟��'^j�������F�:j�Ad�`�r�෿i��	�SY�<�	��	ܟ��kyZc2B�
⬖���9���2xDL��4�?9�(<K���IH,oZ��37�ً|�^�`�n@�M����?���?����J/Ob��O y���<0Lu&�N�]j�h#7�����0���h�S�O�r�]#o��͒eL�9%�����X��7��O����O>����<9���?����~b$@�J,�I�W*�a�E�H��M�N>SbR�X�OLR�'�¥ңh����b$�1�R�����}/�7M�Od�:�F�<Q��?�����Ӷ��3%|f�)��U�Sp���o}2�!E��'���'�r_�@{T�r�vi���*~�h�3�ğ?�D�'��'��|�'�R��3V���X-����&�;��X��'����,�Iğ�'F.���П� b�PHҳV�Fm� �����SC�i��'��|��'��)@lm�d8KJx��J�� �XA�A�=h��I����ןD�'��U##P>U�Ƀ%���ʙ�{QA����pH��Z۴�?qI>���?�挀1�'�6��Sc�	\���2DH
.nc$Q�۴�?����ҍ6^�'�?���b��E��"��c��08��U��FsW�'q��'�����T?I2*��`'
�&6���ak�D�s�(����?1��?��'���P�#��E���P�wB���`� �ib�'��$É��)���<���S�/�E�W/�0���W�"���'���'���Y���Iϟ$�����\\�c_�|��ea���Ms��A��������U����,Y6_2�Qx�I��O��Ul�ǟ �����C� S ���|:���?� �)D����O��*�IJK����'"�Y���������ɍ
�Tl��d߻H̾��ҮI=P����4�?Y��K5&_�����'OɧuGjE� �6�����[�L�����?9/O����O��ļ<	�#Zl&�0�1�,pzT����u!���Q�x2�'�"�'0�̟����Hg&$`�&�]��p;��[�iZR�
�ɟT�'���'	�I���yT�a�s��[	H���
.�m����ʦ���˟��?y���?��U�Y��oڕ�ҝ��,��
q�J�*9�5�x��'��	����O^P��'�ұ��KE�?�,�S�ă�M�׎}��㟰�	���@��p��O�h�C&��\`�a�a��=y�iA�R��Ɉ6� ��Ob�'��\c��p�] x��i *�Y��ZI<����?q� �PD�<�O�0�p���0N�$��Ӂi ���ش��d�9�dAo������O��I�t~ҏм
�\�pM^i��}Â�ۓ�M����?!B+�?����O��s��}��R�:R�B���{N���`�i��%8�'���'B�O�)����A_��2'� 8���c!X<F�v*J�R�9�y���O�}ჃH+�L1�t���4�qa�����韰�I�y�:��M<�'�?	�?���@w�8r��=�ʞ%�p͑��i�R�'�R�P0'�T�g~b�'��j���P��l$<��bꁩC��6M�O�E�2�Yg�i>��󟜖'��gD7 ���#C߾(�RE��fӎ�D�#2b8��<�'�?�*O �D�-2�����'���c2@^! �`(��n�<����?��B�'p'�+q�X��CdP2U���!&�O��5f�Ø'�rR����'�(����P�ђ$C_&�AP�����9m�̟���T���?��,��-R�YƦ�A�.PvI��Cϑ5e�����(�D�OBʓ�?�vnI���	�OZ�I� p!B0+�?�"�Xs"Φ��?A��?����g�i%�`�1f?l��dj��'�EI&�p�j�$�ON˓���X��t�'��\c�Z�c�Ŕ4�.!hg� �^Z��۴��$�Oz�DH�J��/���kL��TL����G�v������̟9$�\��P�	˟����?���u׮.7�E��>d�\లA���M���?YdHՇc����<�~0!B#v���K�G�D!�����u�V�]�L�	���I�?і��	B�<�rM��C�6�d|�$�V�\�@�nZ�x|N��'�)�)�'�?�4��8?H�C��=n��P4���5D"�O����O\4pD��_�i>��������)�'M�u�����0�Z#��M���?Y�d��Q� X?�	�<�	ҟxҴ�ç K�Xӵ!Z�)��%Є��M��9�m��x�O3��'剧 �5���/S�9��ZN8a�4�?����$�?y+O����O��ĭ<�S�	�gt&(( NX99n 
ЊYM[`�qW���'�BR���	�����?F�
q��L&5	PmH4�IP)P����{�D��Ɵ<�I���	dy"�U����9�K�y��)�!�=(`�6M�<�����d�Op�d�OX��gU?��� 9~��58#�Q�X��+f�f���O���O`�7�Q�X?�����<i�.U�G-F���6u�ԕ�ش�?,O����Ot��ߖJZ�d�<�!�5^����N�{�c��ԗ#���'{�S���������O����X���kSh�����jx�CfOJ}�'�B�'i�@Ο�ItJ��_�3�F98p�<m~t䲐O�Ʀ��'�X��3IwӤ���OD�$���֧u�+I7&h4I�#�q��A��β�M���?aoJ�<I�Q?��_ܧ<�> �@��{B��@�.���l�$O`��ٴ�?9��?1��*7��kyr�t��TC>�>41Do���6M�.��0��.�����cf�v.|$0���,

b��P��M+���?��*��5J��iDr�'�R�'�Zw�8�p��q���WAӖ+����4�?�/O�T!�2O�ӟ@�	����N�>eW
ll�A'M�
�M��V�jvQ���'w�]���i��a�+D�%+�Kc��&|Ѽi`��>�Q�G�<����?9��?����D�?l����4�F���1�(`�L�*U+Ez}b_���Nyr�'pb�'�T�����E�LI��@��BH�A��3�y�\���	П4��sy"�߻�8��h�D�[=�@��m�j�Չ���'�bZ���IΟ��I�h�i����� Ҙ:��.XL���GpӤ��OX���O��d�Oz���(���5�I۟l��!��]����V�Q�B�8�f@��M����?�����D�O�� B�7�ɞ9�@`CA7�Z(JJZ�)��g����O
�d�Oh�!p#�צU��ß �	�?��
� �\)��ݲlD��*��A�?u ��E�ibR���	�DT��SH�i>7�T�k|n$���ߴ��X{�d�w��f�'r���n�6��O��D�O���������~\�#�7��<��@A��' b)�#3�'=�X>M��x�"�ì]����W�~�P��i�$��%������OB���4��'��	&,�ypH��JF���5����Ubش}�y̓�?!*O��?��	���q����i����+����4�?a���?��Ί�@��6�'�B�'?��uw��A�,��#���[׮�!�MK��?��P���S���'�r�'q��!	 <�!��f��r An�6�S�Ά��'�I��@�'Zc;ֈ��:v�⅏��T�P�OV��':OB˓�?����?-O,,Ȓ�D� 		E��T9�X8�c�7����'B�؟4�'C��'c¨ƶQ�U����|�p0�Ü96F�қ'��֟���ؖ'׆9��t>���T�.�<<�FI�i� ���lf� ʓ�?!/O"���O���̖U���)7���A�M[�6L	d
ּ2��lݟ��	ğ���Uy��΄ꧯ?�c�G�(P����.�����X��f�'��Iϟ���џp�iw���	K?�E/ύ�H@� ���d�8�f�A��1��ٟ��'�n0���~j���?���47��#���8YX@� ��o�0��R���I�x�	Z����]�W�e��&e����G�xG�}ʁ����ٗ'�v9j��s����O����&}֧u�g�:Y,���k�~�h4�MK���?! o��<��]?���Y�'x醥��m��Ks'V�b�P�n��;E�aAڴ�?����?��'PK�Ily�/U�-=^e�g�ڜ��$���x=|7�S)#���<����O2�8G)�ة�B+
��C".��DB~7�O�D�Ol<�1Ho}X�\�Ij?Q�AM�+2�t!�"I �[c�r}�Q���.?�'�?Q���?Y���u`�J��	�bq6�r�	�����'��Ȱ�C�>�(O8�ĥ<���릇��U�<�@�,z.T�`��L}����y2�'���'�R>�	4&��@�曆X*,���a�2Ƕ��`�:���<�������O����O �Z�H���xҡ�NR�r���
b��d�<���?����07#���'D<H���ҿ6�XH��I1V
�'�"�']�'�2�'���B�'
�y��.���Q�F�
&���p��>����?�����Lژm&>��D�ܺ8׾�٥,X3���0M��MS����?Y�h��IΓ��kD]B���b�c�D"u�նiw�'�I�Af��rL|������(Ȧ/6��*r��g,��2SηQ�'�r�'�b��'Cɧ���v~R�x7��=1����C9(A��^����E]��M�T?����?u�O����8Wݪ}Q�ϟ�~>P���iC��'������'pɧ�O�����ǂW:��f��}��ش71�q0պi�2�'2�O^\O��Dܷ^���[u��Wp�z�Q�m�D�o�� r�?���t�'���'W�+�(EB��ΰ_5<p!��'yr�'L�4W��O���O��I@I
�3�#��8����X�7�)����.��?�������	�B�&t@G
=$׸�ϑ%i��4�?�`j�V�O��d"���x9���F)�"�13$��Wɜ�pQ��Ӕ�j���'�b�'?�Z�P��1��@�ポ�{.��
��`K<Y���?AN>Q��?��o	;���E�@.�l����(�y����O$��Oz˓V��˵0��D1�OW���u�D�]����_�p�����&�t�����ڥ�}���͆o]|��B�ʹM�4(�-���d�O����O�ʓ0��}y���Ǜ�;�.�����F&j)�׌$L�X7��O�O����OZ�����O��'��+�!��~J�%��a�4d/�q��4�?������F�6$>E���?�+���v( x��ͽ�^e1V����?����l����S��c��n�[S�^�cp�q�
�M�(O��Ig�^Ӧ0�������8�'$X+"��\^R,��I��+|(�ڴ�?q�]��D���S�Qy���.�"�(ђQH�;xBf�n�
q���������	�?�aM<���$�,�(��$"H�;DE�=�\���ib.�*T�'�ɧ�,�d�27�d��eI֦3�0�/�|�^@n���IӟX�ݵ�ē�?!���~�ȪE���E�ݣ��*#�2�McM>A�O�"e�O�"�'��jQ�2�����_�X\iz
H�N�$6�O򀳱�_k��?aO>�1>�f鈄��A��XG�VQ8	�'ɦW
]�	����֟Ж'�J�J��2	.\�:Bѩ=z8؂E C��b���I~��ޟ����j�R�r�jEU���/�p�,d7�w�x�' ��'��Q���7�C���Th^�*<�.��I�| �ɞ8���\6m�O0�O��D�O�)�(�OdT���I!�XH3���b��
�O�j}b�'�'���'� ��q����O�ԱG!��l�y��gp��Y�a�����qy��'��b�O���O\�jtⅼ.�@:#�O�PyxE�e�i�B�'f�'<PM�U�dӸ���OP�����	N�I8# �zd��+d���`�m����'m�Ȅ����'��i>7T?B��۲dG0 h��[iC�v�'?r��ܘ6M�O���O&��䟖�$�t�(q$���F� ]2f�"|2�'M�*�*��'S2\>���ThiFědOpA�@.�>/�tHr�i�ft)C�i����O����	�O@��O,�� T��ƕ� cx\"�n�A#�x��i;Ty��'bɧ���d�'��8��C�D팑�D� :P�T�`�lӂ���O~��^
u��m�L�I�T�����]����s4E�z%ȉ@PCF�ZL7��O���)����?��|�)[��:G������Qy�E�i���W ��7m�O�D�O����D�O��(f��:qFDP��;n�Hc�U�`h��g�������Ißd�I\y�)�� H�c�y�3�K�[��T��î>�+O����<����?a��\(�#b���3h�!�u�؇;i8t����<q��?���?�����ǎ1W��lZkp~ 9T��V#��[R��!�М;ܴ�?����?���?*O�dL`C��ȡtU�4�0l�K}V̐##F�K�ޔmҟ��	ߟ0��[y�Ѻ;�`�'�?I��Ձk�<�1W��'�=�sEIV�f�'���ݟ����`
u�#?�禱�X�q3��*�ɛ#J�x���kc�����O:�#I�Pv\?Y�������bx��be���T/��8&U�	m�T�O����O���X�*��$�O\����B\D��hE��7pֺl��͏��M�)O��Xu�֦��	̟����?qڪO�.�P�L�����/m $�>W���'����y��|��I�
i*St�-=fƬ�pm�3*�����e:h7��O2���O��I�m}Q��HcM�`$�s���SB�q;�(E��MK��<���d-����0�(١�A5P�W]ą�1�D�M���?����|��7S�@�'T"�O&��t"U�+�6���Ϙ�
�:��@�i��'���X�����O����O<��q���<���H
�#:��jR��Ħ��ɟ{���O,��?�-O.�����K�c�<�p+̚l�l�ix"���y�'a2�'���'��I^6<AJ
Bi zI�/�
Sհ�ѐ���$�<������OV�d�OjeRc�*_#���@��]�
`��G[�9*�$�O���O���O�˓`�JБ�0���85�6X���*c/�a�2U�i��	����'��''�����`��ҁ����������4��6�' ��'4�V���5�̶��i�O�ze�'_("�a"Y�Rh��'�F�E��@yR�'4�'(�X��Ol�ia5O�F�zT{WGۆO ��f�|�H�d�O��<�z-ېU?���ӟp��8-�}��-Υrή�*1M%~��%ѮO,�D�O*�DI.|��D2�?)��ɒ��Љ��)ǄL�x2�jx�<�2k�L�i�R�'��O��Ӻ��Ϟ�)N�q�gAC-�Zt��aX�������Q�|�'�d�}�gk���HM`w�Y�&��@�W�覕B@%��Mc��?I���7Q���'`�$j�t����玉v/~ap�gf�H8��9O����O��d4��П�d@��2�Տλ5|Py(o��M���?q�]��c�Q��'���O��G,D_y��)1�ٙve�� "�i��[���dem��?�����LK"��&ᖆ`�D�s%��M�+���'\���'7_���i�u���ͳl�H`���6)�X�cd�>���]��?y��?A)O4𰴮�.v&�$��ό@�|�8C��t�Z��'m�	՟��'l��'Ur���e�@�P�վ@2c��,��|��O���O��D�OʓDl�YS7���:���>=�����+x3��s�i��I埌�'���'��O͛�y�Nɜ"i`@`U��b?.$���]����?9���?�,O�@+��E��'h`H�v ��}��0��� �;��y�үu�����<���?9�*$�̓�?��z���oK4}z�@8q���Ӱi���'&�	�i�dԙ��\���OH��<
<�)�M1`>�;6�	 J:���'��'O�C�.�ybQ>��p��c��YO �c�[/2�ʁ�P#�˦	�'P�d�Ue|��D�O"���Z�קu���;-��H�g�Y(+D�@7�*�Ms���?�'Ou~�^�h�}��f�-�N�����tL)+e �ŦY��������蟨���?E�'���[��@Q�[�,��MR��C�n�~i�Ot�r#�)�ޟ�Q�&Ƿ!� r�E &f[�e3Q �5�M3���?���n�8�rq�x�O���'��l�@V�&����i;E�� ��"��'[5"b�d�����I Y7��ᮚ�@��ʵ+�&'�Aٴ�?q��� ��DJ���'��'�ld�T��EbvE������$���g�������I۟��'��A��GM�8�aEŅ�(��`����+X�vb���Iퟤ�'��3O��8QcƠ>lܳ��^�GH�hH ƚ3��'5��ِ�/E���E�x��ȳ��ϙ��	I�4�v��E�ۧ�Z��3DE �!�d�N2:��DY|�Ĵ@��*#�qO(0V�Րgl@P�aA= �b�k'Oiaf}�� Gp��B�[�Oo̬[�m�4;u`�Y����&���4GοɎ�Ґ�Ȁo�y���V�{<L�Sj�*�|6����|��!Ί�w�*u�cAI��Y�"MU������S<n����	��!��M�A�ȡ1 ��3v�-!�'$j��o*�I@��,�6�s@�'���QN��ps��O�!U���B��USf�����3/v��:��l����K/j�R0d��ǌm�� �Îb��vcj�I�;��ӎ7t�Z��3
�	�"I��t��'�+��?I����OНy7e�w�F��A͐�a�4l�@"OZ�˅dځ $=!fF�n>&��',�#=qւ��: TY`�AA��@��e,�f�'5��'p�б���'��'���y�o��b�\�S򥈃'�h��sƗ=��)A
Xa}"���>=���L>��B��Щ�� QR�(�����<+��c*�>�UO��0l��>�O� �p U/�
W��1C��<��y�7�O�D�Oh$��/�Oq��	П�rb	T��T�����:��oh<�e�VHx��v�A�����
\~=ғ��<QGJI �Q3��w��H��,џB���A���?��?�����n�O^��e>ei�芃�<=�ԁ���6��_�jB�I�'�zx����
VR��-��0L~���+�|��f��&�z��V�"?��p����<ɂ�$�Ox���O������P�I�	�a�=l��	q-�"�!�DC,bPĠx$c�+2�<��iڢx�1O��'�削U�$��O �䕗__LqA0aϷ��Gh�(,� ���O	�� �O��|>18s�\�+l}��LQ���l�nIq����Iy��+��77ѐ����s�]`'h� ���MsH2L�ɢ%]	$�|-#�l8��)1��O��$�<Ѧ-ݣ%@�Y�O��)8�) ��Gj̓��=�1,ϲ	�6]I��о:���K�
<Ƴi�H�b�Ö�4�v��c%w�8�' �I�e�N��O8���|��G;�?����f�dT��WEh"��4�?a��IU49��̈Ċlj�G�a�*���'f�jњ��{��X�5� �ͦO�E���d.�ۗ�W�n�"}�� ��	�2�S ��|�> C.�B��8���'a�>A���x�r$CchP R�T�eg6�C�	E�h+t��L���
w�3U?���^�'b�db�jW:5>x �0t���2Fl�P���O��Ĉ�5B��g�O@��O��4��͸%g�+����΍� ���%>�	)c����'�b���$�xFd��CC�
��I3�{�K�k�nх�	�k�^���U �G�\�>�����\~φ9�?�}�����I�d���kjX�;�*�`�w~�U�ƓLW��kۙv�~e���D�?o���'�"=�O8��,�J왖! !�C$fX=NL!RH�)e"����0��ԟ�^w:b�'���B��ݲƀ�>"�F���+��	c\�!��%Jc6���ܿ}�$T��/B�m����)�1cB���L?�̤����[�@��?f\���-�X����]�!h�b�'R�'��V����v��P��퐍y^�ٱGI���x�V"OЁq0�U�GSF-{�KǝSľ��b}"V���$��M���?��,� :�aqIS�6/��zA�ƴ�?!�B�
��?)�O���@�'ԤIظ3H�)&��J��5_����o�(v����"��t8����@֦m�3w�Ƒ�@m2g�ӌB����č'�&��B�5B��x�g[��?���?���R�Ȝi!M�9�e�K�c���j-O���%�)§�r���Z�^3�][-��r�Ն�dK�&k-��=��̏^��@F�Ͻ�yr[��������O�ʧ0a6��!�̉���YB�a�`�,�������?%�قr`����	�>Of̑��"bg�}q曟��i4U-V0�����anJ'O�('�~*xiwHZbn�H�R�ؤ�Q'H�v��'X'���eʥZ��pתC�L
ŧO>䃑�'�"�ퟠ�i�n�,P�g��\�Έ1� 1D�|HQ�E8��}�����L�E�$O<Gz"ˎ�FEĤq��58���^�	����?a�"�40�/ӡ�?���?��Ӽ�b	5M ʖHJc�~�(6"ϡZG�p�7�L�[��˛�[F�Ҏ�L>1eާ'Ą�Y'AZI+��P2�d�]SQ�U�Bu�G�FP1�}&�����L����L��[o�;bC
՟��	˟|��L��>˓�?)�G�,g� �E�G�>�G��9��x���ls�1��,?�ղ"M�����M�'I�UyB�Ěmt�@�OݩH1��!ч�:e����g�Q��'R�'iv�'�?A�O���%.�NxT�Y3"��_֢-�U�\	d��B�,��M�Pǐ�ul$��M�oߠ`�Ο,<LiĤ8f2����?Y��!r�F�]�.�зND e,}#g�'�2�'��V����W��\�R��)� �1�KQ�}
*��ȓ8�8�T��,*�ĉ!���l���<QZ��'�@��/tӰ�$�O���lJ8t@B ��ٱ|�^��j�O����[��D�O�S�D'��˲�U�l�����'�6T��%�]���I"H�0Mw�l�	Ǔj&��� I;F�Y���O����N��B����^�P���p<�D���$�I���I���R�_��@h��]�N��9
V��<9�����*x��K��8�btrt/�/�>Xp2OԅnZ%^�!�dܑ-z�M9�i�$1>�Fy�G�6�O��ī|uEK%�?2��"�qa���c�5��,�#�?)�~��pb�'՟��[!n]�%t*�jʧ*�� ���@8�{����1����O��D�\(8c�y;C̄6v.#}b���~�4]�%[8/Hd��d�Y�ʶpQ2�'R�O �π  1�A�&9\Erqlڤ\�����$�O���dF;\/l�	dOM2�4b$�ъ4Hax�l2�RS*p4FV >��K���6��%�i���'�" ��!x��r0�'p��'�w���q���CCT����2/y� (�9.��ɯ^0Ƙc%c>�3�$�:�(�3���7��Rx��@�@����3�,� �C%�3��\�om��4��"��}���m�p�mڷ�Mk��g�6A��S�gy��'�jlX6�ڇt�j-�d�>k&�[dO��<1a`��`��w�^�xw��<ۈ���~BR�00'�\�n��	ӳK�:|�t!k@������+�������	��	�O��Su���2�W�$���ោ-�.}{g�h��̋��=��m��B�{�(p�&u�y��ɇ=��I0�T�j���S�5J��\�^���'EB�'L�ǟ��?a��ߛe��i��OYˆ@ �`�k�<��*���A~iJE�c`�`�	���hy򊂟.7��O���M+1���dUR*Z��∘��D�ON�x"�O���d>��CH�P ���ŀ%g�(oZ$���+&ʉ�Q�b)ۥ,,$m ����0F�T����R��om��mb��1��Daf�� ""�3B�'�¼K��?�(O
�a�X�8�� `����>O|���O��"|�+ʼ=�hB0,R*8�8H;J|<�i�����E�J9hdH1����'�ў"~Җ猀w� �#ÞT��ݡ�� x�<1�ԋDx��*�
�%i2lI��p�<iፒ�p!��"'˕ukdm3D�i�<��k�7 �SUƘ�<1�B�Jg�<����+Ȏ<�Щ��t������^�<a�M�[?JH��X<��7m�T�<��䏋sW��!Ꚃ#ʨ�q!�P�<�p�C�|�\q3�Ԁ@�R͈G$Ht�<3��0eAs�%�9R+N�Y�u�<	��~J�pK��J�xk�Iy� t�<y���2i��l�B������^q�<���(e����4��P8U�E�<���9��`��F�8��,�B�<y'E6�@�Y�hJ�+&��3#�}�<9�(Cc�L$C�ʅ��HhUd�z�<Y��ؖ8k���͓/����u�<��ھp�X7��h;�)�'
U|�<Y��	��m���G	2�k��^P�<�V�  �JL�I	Yht�e�M�<ٰ�XU�0�2N�9F��ŢQ�M�<�q
D)z��HP��^�[iRH��a�<���ߗ;f��yAdW�R��`_\�<)�%��PvB���.��Wp�i��*\�<���to&HY�P��P!���\B�<��'��88<�a���*	Ʈ]3�Q}�<��	^�Ur��V�/;��}��+�A�<A@h��U��]yr���Z��u�<�H�d|
)����jw���D�Tm�<�W)ۡU*j]AE��n��)yp��;�X���5�� �I��Gǈ@�}�H<Eg��	�m-@��t��_< U9%������it�H���� @:�9QVi\�0�ع�BϞ9k(	 �k)O�}1��;x"�qX��F�Z[(<q�l�7#H`��#*�U�nu����3�p<��8KN�tb�j�X�r��˝�Y����,[V*�i��ɫ<Tr����d�ڬ����(�~����<�r�*��6ل�0��$q�� �&lO&�� &�;D���JQ�N��Ȱ!�Ҙ"���bҨO�;����/�::��'FuI�O�*�+���f�u�7�[�x��r�I�D�u����0$lb�`�B�X�����TZ��-�"/B��'��*�c��:��%H��p8l��剎�F7����Y� � ��F���hpk��~H��?Y�#��gOV�'�(O\$1 Hߤ�R�y�l��=2|����U2C�'st�B�阩`��ۜ'��V�C3?lq �̄��%�V�\0-�<3���6G����ėbU2e��K(!n�ԈȺ6T|�'�Bҩ �1��rì+ڧjsru��B�M{xS���O�$�!��^}� B�:r�rt0�#���rjȃ��y`�4+�!sV`ڲ����#��ӷ�:� �#o�a�1r��Გ� �mbp0�5��5�65Ey�fB16d���q��D�ʺ2��a�'� ����NԌeMXe��GZZ�¹�!�>O`T�R�D�o�Ԣ�&�;^2��� NՎaEHE��{@ΒB�ҌFmY-u:y��d��k #��y���~���BH޲8ҍ�eHq2Y�3�*�yBd�u���J0E�:.^v�J��TO�F�S���D����mK�����	�7�^EJD�X�X�*�y�"�	{z�:��T�@��ʑ�S��r��#8?i#FE��$
�e�1mR /����z5�|�O�3���̓�|�	���d����]Wr]H�I݅*�\�'����,��iZQ,S,Ԟ���C�H�>p�5�ce�bp �J��e�+�HOL٢`k��<9�^G��A�6ƅN>&}jv�1!�e�w
A<3��#�b���R��O$?/ �1�Ѐ���*�
5)�E��
0�I�~)� ��'�;E?t��c��&i\c���k��f�\T�J�~���pK�+e��X(�d��Y��9��=��B����P�CԹuʜe��
��j��'������Z�y&~�S��]��hB �?)���c��q}���q��$P	����O�@1�S>Iki ���Um�"�֘����Q�<q��ӆ^X��҃�D&#���d�.�p<�GC�S��!�G��p؄��3yj\Lc$J�!p]d��a	���=1 ��,[�,�D'r�$�&B�<���f
�3���R��>9u��4����H�<�4�|2-,pR�hC���(�L�y�.��O>n� *O��0��m�T}�uC1iδ �c����O<ɗ�CҘ�sp%ŗaޤ���-س<��ї'߆�OHa��ѵԸ'|"�b!o�1/0.� �Β�.�8�	�/�Vr���<���w�2�s@D�#O�����/�85RP�On��O���O)��i�#*:�5(g쓔��w���R/����'��r0o �s�ʓF� y%�ǥi��а'��5-vz ����a�.L�A����h���� ���.!N�V	�!/�\�2���5c� �@,O�!p�Ü�OW��' ��O�	�N��� ?h5l`-X�U�2��N�P�R��6@V�TZQ�������'��Y�獄 ':t
��Œ�B�k4�nӼ���'A4�ZN�擮@qO���5��?|����
�[ܪ,�Gj)�����	M,�8�ǩ�r�����sf��|��dF	�❢ �>M&rA��B�DF<L倌�¸�MB6���a%6Yb��_�{|�yK�J-Ld:�Tf;?��'XHu�/�*��G�O�����'�E��*�v0�B���}y���G�	bL"�q�W.{b��W�ڞ|����On�� ���{�.ʂ4$8�1�.�h2�����gi�-�7�`D�I42Z�ҧ�t�Ә��x%'�c�45�Ǥ���MwꅞQ/�e�f���Fq�U����ǟ�I^�Ozhi�QU?9A�l�Ls�ɪ����W��y����?����O�4�4[�{�b��j>"�v'�!�����?�y��+�O�ULX�Y���n�����Z̕O��0˃��t�,9�q�՟N�b�`���XpT�Ћ��A�M�vL��_!Ʃ�B! �D#���T�����D��OH!�C#�øO�٣������if�ֲ3&�������ArIVu�'K͚ �J�+�HM��U���@4c},p��H��Q��a����@0��
7�T(�O@H�d��O��R4�C3Ҁ��۟����k�Lě�႒+t2�CsX�\yb*ΤL��\��	��섁�
څ�rl�vM�%Z�@�:�'IN�)gJ�+�¡�S�J�k{<�B��"�ź�|e�U����d�N��'aP�tR���)rɓvG�7;�v�UF�a%hy
�*�	7T\��l� ;%�tT�~�ȑrG�{v����-��̎��xs@�&o)��)ˢ^O�y�T�G��i�
��ywl_)p�qY�n଺��ǽQvD� #��~c݇`�~�9�':�i������'ҺX�eΆ.`��t떉�9(-�[#O:Y���C���c�\�rW��zË�	~z"�ٍ�L�(q��M?�� �3�?�b�O���g
�?��F	� '��A���!7�IV�9�;AȊ%��U
x�9��I89掸��P�*�d"�
h@2ɋ�5��<i�BόmO�'��ɖg�8{SH�	�̬�=�%�$��jp�ԁ}fd��̏>��CV�P�f���aJ�P�|��)u��ht�ġ=�d���3֫I0O�	���<r�7o
*�MK�Y{����O_��p=i5mS)���H�.�2p5�a;v�߄v���3"�s�Z�Z��%L���J?�����Rjۤ��)��mHvb�s�I�
.S1�G1��� K�iK	`�C�'a����G��,:�16���0���TP�}0�)Ƞ�>�%��2�p��I�sFf�R��[� h'E��]QR����I�M��՘'�K�E��Ҥ��'��%E�x��7EH�DT�D�]�(�ɑ��T��xS�ӧ[Ҩx:��\�(�
E��0|�!���SI(�o')�����Q��ͺ0 ��k ✸K�z !�ʌK#@����f�N���[��Aئb~��O��u� H��vk�ѵ%��4�&䩰�I'I �y�	YS��� �:�oƙ#< Q�@�;�b���HyyB�
!8dn������'�n���Ϗ@%P��2��25��C�Jȫy���)$�'���c!�Ŝ,�����J,T["��6@iHmh��2$(0��J����pRd��"϶ HGbSe�� �D���p� �u�L���K����"�2�	/���&��+��AYc�\1|��c�� ���<}�~�����Ƭ�R4��O��ѓ���N��e�J#�"��I![Ԅ
B��$Ka8��]M���qH]�`�I����^{���҄`-�5�uO>�@�^(e[ L
�*O#�0=�B'���ywc�X�
�OG�<�ϊ��?��H1V�{��U;dl��#b�|�N�:u�ɉ+�<K�vd���O$'V�qx\y���=9Ǯ�Aѹ( ��υ.@��%��[Ǵ��;r�@�H
�DEߟ� T������%i�J��U3��i�� kS�y<$�U�F�*�ة����ot�hp�V�jir� 8�BI֩BO�G��тw����3�2*�j�A�L�Q��Ոc
�gUN(�V��8�p<�R+�	\�T;�'�ǪS?y0�l�N�� o�YD��1,:�у�ڄ��O�z'��¼CP�ʻ�aC�=1d�8Qu��{�g*�<1"�O�3�*Y{#nA�7Լ���^�8���i�M]+�HOZ�ڢh�:�{E�ŝJ�<���*�Z}���
B2d��ؓ�DY��H!�(���J'a�����Y����xt�v�Q�VI ��h�FA!�Q���)���"M_(��%�ѣy
4p�(� ��OP� 6``�J��B�B5ā4�i$������i�Q*P��0��]w�� a���8c����ϓ$]A^R��"�.�1�C�ɟH����G��B���eD�h��ܲa���6��LA�$��F���b�o�'���alz�$���AK�Io,��NO�\��O,�IS�굑W,և(�R-R�[�T�0�i��6��8�2����HO���%#/*j�ʰFT;��@���3עW�b��D� �ޏ+Ϡ��}���h��Æ�L�͊$ Œ����0Sv�
��$�83Rj|�` ���s�
��8��+1�l�S�'���0mG� �>����KKz��%J��F�$x���C���,��
"yj D�7���l�E�'7Е��GH0%����D�(�<e���d�-4%t��O�	�������GAȠ��/�.* 3�����^$Yaz��W;��hA��9�0U.!��3�h���"v��**2��q&`�O�J�7͘�X.����'6�rf��*��A�C�Cax�)�;p[��OZ9Jt�Š9�8�h�#�B�rLSN $,H-�s��f�b�#� �$qU�@ƂՀy/8�=	�c��\��y(S� �G��L?)`�S�,8��z7f��ݴ�(O�Ҭ�"U�~�9!���A@��B��mM�(1��W�(y��.d��C$�R�^u*���tb��pE�[R�X̓J͢�8�����D4�ԙ�H��J�#�c�O����5� ���8�
O�5�r� ��� ؐ1�$c� ��<Yg�A W�2�Z�M9�:�ߑp��e0�n��#�BG �[T8">9�C�L&��vh�h��r������̹<�@18��
9O#�<�q$}r��52F�{���b�>�;����'?L��*�84s���"煄h���'*B�A7��o�^I���A�?�L���D�jT������v��,����7Ĵx�B�8� �h#��b؞`R�c?N���d�0p2�ED5����d/�OY{D�H#g�&��KV�q#ֹ8"�8�O�� b��c���K��-���@�&72b�
ϓm��B�.r��
�&�1/2E�c,�(4VI{tJ��cfR�s�G+�<8���s��8`�!�<2�B���'��\���L�t��($����D�04+�)"%�
�"!J�5��!�bY8B�_:�6�q��[�8��b��s��K�x ��U"��c$�T��c#� f�r}�T*�U����\�C+�b� �%��Za���Q)�z��&�2�*�b[�L�&e�.7}\�b#����J���
��<a���
04i�3M�0?�lB$$�yҎҟb���J��ϲ~l������<I��ߒ>�����=Fm(�+��ׯMҐ�r��6V�p���0=�E�_;k�@9��b&]?~l �@�,|kT��..t2�0��^�	P�2�2��>�d���N�?l�p�у�yN�)ԁ��Pd�8��)扜V�d�:���[�h������8c�����]\�� );䈪T���(��k��8K"в��'�����ǀ&��Z��1��`O	H��c�!�u@��z��h��׊����"DL=z��ԙ�'� ,""�	:ހaK��<�F`2�'h4y�%I�74���P8H�Y��+�m�"�Pk�l ��A�;�OAA4�<߬Q�Y ��u�F�	|�����Hl ���%�_/z��@'�.Z����~���q�V�I��⟴�V�P�qUÿb���zԂ7�J�(�"l,�����?EVD���Q� �F��Xd�bcϧ%[�K��--pI�aH�e��]6�'m�����,5@M�&^�a�X��NP���)�R�.r���5����
���?��O�%��y�QN`��H��#u�����0bE@!�5D�x��Z5?L<{���~��8!Á'X�T��ű#F��D��:X�e�K7�\9f��>
�9	%�q�Y�n�~9X���ط V`��'/�O��uO+���Ñ�w��"�Z˦�Y�E� X�13se: ���d��%��	���17o��&�d�3`J\�����.L��a�H����x�6o;0,`��A.���2>�N�x�`��"���q�JO�B���wOx��@�q�&l�S�כAP��`"O�X������Z����N�\�=��"O�EcT��|Ld���a�.z���"O�����M�T�S%ρ�3����W"O\e�T�ٸ6���ЬAL�Bl�"OJY ��^,����͉h��r"O� ��`��J�"���C�KJ4jr �C"OR<�0��mfF���I,	p8�i%"O����3	��#��b[����"OR�J$Y�QW�	�<��i� "O�!Z5���3� ly5���%��%��"O�#5MO�]b�\�$�mC���%"O���4��5�T�D_� :��"O��ZU�� lF�QÊ��(dL:�"O
pu�̞u���s�E���ep�"O	��^��9f�ǏU��� "O�qD�I�a/���7A:�@�b�"O8����֯!�°��m��CR"O�� N4A2 kS�[/� Y(R"O� �eO�.���)��;���"O��+�-R����e��~�:!"O�Lh��L�T=� h�MC�8ɰRQ"O2��Ã
{�%	��Έ/g�T��"O��h\�[��jgMZ>d)�"Ox`�L�:�Nl24�@7}E��"O��k�aE�XNv-A��ʅ�.-��"Of�:�d�-o�H�0@S�V�Jp"OL(�D/���6���̃ �Iے"O6̃Ǯ�%SْmȣF��rh:G"O���'�!d,����=)���)a"O�)&�~d����+~�e��"OV�"��Bb^>d�)3
����"O�Ҁ]�H��䒗'�)�ܜ��"OnH��E%���+��E [��"O|9�ňپJ�d����3w<l���"Oܨxa�@�~ܸ��LU�'-P ��"O��.G(cڜ�3ClPk"�Ī�"OfL�����Y����K�o��
&"O���F��K>�YCJ3.ސSV"O��B�&ԟ|u��˅h�D�qS"O�p!�g����0�D{9N���"O�,b��2]���?0\)%"OJ�� �;\�\ ����\�ސ�r"O�sj�l�@@s����t�{F"O��!GI�r��yX���-��U��"Op�{�5+�x<��˟D�Zi��"OD��"OaI�X� X)ò���"O(\�1 �%��CF��+�<�)�"O��0T��VJ�{$��p�&"O	����t�xɣ�)B-

�:�"OezUr�R��F��$Ty�"Orh�wdS�Zu�=�t+O���6"O\|3�J��^֤��Ɍ-$�� �"O�qbЀY��*찤�Y�Jl&Y�P"OV��f�տ�01Z���sd��@"O�-q��!PԌ��V�E�Z �x"Or4�M��E�p 9d
 ?�I[�"O^���J�/x�M�������q"O���6E�<����Q>mҍ�"O$р�H���)Vē�I���v"O\$�!�ڇj�d�V������E"O��s6���g�d��*�R"O(`����.Dd0k�!�l���"O�S�̏�oƮ�v :Al�q�"O��#�A�x�)��	ݹjn����"O8�O �q�q�I�H\q�"O����g�p9�
�$zX8E�'����Q� *6���f�ҹ���d-D��s ?��l�g盪O�E�G)D� ��j+g��@cd"�8:�l����'D�� za��	k�I��`��YS�"O�PiReZ6��M�C��bb� �"O�4Qe��vY�$K�J�"O�l	���_p�f7�0s"O��s�O���d�{�O_;N�9 C�$!\O2)��Z4.H��K�G;p��D"O���J�I.*L*%�}��5��y"n�zj�y�� Z�nd��.
�y�ðl��x1�5wPasdŜ�y��	�(����O,�@�q�ѽ�y�]?U2>��5)��I�U��y"��I
,�cb.P�/��(˕Ɏ	�y��O�b<#��]�q�|�Bu���(O֣=�O�:ai���8�P<���.��),D�d*q�c�IZ 4ض�Y��6	r
�'x�dq�_�zr�IV�
��P�	�'���s$	��=��cU��R��'��=������Z�i��1R�!��'�@H6�J=��:ЌN�.C쥹�'����DD(Kxa�fON�-�Q��'�u����"t9>]q��®$����Op�=E���W�aa�d!
�(Nlܠ�J�8�y���@��:�O8z�
q���yR�,W0A�G']���ᇥƎ�yHR�x|��qv�i��i�[��yb`+e��E���X$g��atK��y�nvg0A�4k��//l�C$dF�y�I;:�v ���#�x����yB���Q4��DΚ�+��rf�
�y����J�]�b��Ӭ	��ܔ�yrE�r�R%��,���ӆF��y�����b�+��*�J� �W��y��Y�"�V��::��AS�MX��y���E
p��cޤ�5�Xk��B��I�����չW��T�!A���nB�I��x+*n�n��&��f��C�Ɏ*^BI�-I�^�PK�AS<qR�C�9L[�DH�&4{�8�
��O)'$�C�	/D9��N:|�
���C�# B�ɟ"���K���,���8�f��x�C�ɕ戕�Q�[�2��ుo�
&݆B䉸y�U[��i^�0�e�jM�C�I�U�h䚵��+8����.͵�@C��4��d-��N�|��s@�7��C�ID�*d�Ʉ�AĤ���
H5M̠C�Ɉ\'�%�f(5t-+�mDsƈC�ɛ6��@�r���i4�a�"l0�B�I�<b8q�cǛ��(��s�@-?�XB�I�XO���O����Z��ޡdgLB�	/�,�J��1	+P�m�_
������0A�%�2�)�:q:�5&�.D����	6[v����E8<�~Zfk:�Ox�PCf��tć7]�Ԕ���t�ִ�ȓ���	$�a��E���M<��I�+C:t�EpԢ�$�dхȓ"쪵������c��l�v�Exr�'BQ�wgK�6���A�{��!
�'�$�h0� c�mk�K��w��l��']�t��̑�@�a8'��$�Hyr�'�P{�)Q�s6^�C��P0'~�DY�'"����N(`�lHu��솬J�'O|�k�
�70X� 4k?hʕY�'�nD񷩊tD��K���}	�vO��*C�A��udH�
��a��"O�  �
/���'N=+�I�q"O���.�#r�`����M�J��"O�]��@�:AZ��$_#u���8"O��ԀV�g�*`�
Z����"O<dYv���d�Ë/]��u'"O�}�EL��(���Q%Q�k�z٪�"O(H�ӭ�~��s�܈)h�0�"O�ܐ�ב@|��G&��b�"O��b�#��<X仓,YD+z�Ѳ"O���2����T)����4��"O~y��F�=p��P',$���"O�����>E�X�暿R�	#"O��0D�m\�@p�N T�ޥ;�"O�*�,�Kn�m���G�.�*8�2"O� �<;�Ա���x��E�"O�]��쒛v�q�� ���"O
�ZÎ�W.J1ڕҟ4�ȋQ"O>��A�ʻ(�NI96N�N��L��"OT$ �j��2��#ߣ;��Dх"O�}!��#%�Q���'��r�"O��)��-��0!�$��y�"O�uhRj���%x�`E����"Ovh�Z�d��M�@����A�c"O>t�#�`�<��,J�]v
��"O����Wm�0��C+�1Bs�x �"O(EAՃ����A�Q'ݩ
����"O�E�m�)�J� GBm�P�"�"O0���txv��T�G"&0 �w�'�Q�и�F7 /v�+7H��?+����4D�l�u��-��qGɇ3�0I��=D�\yw�,�*�](eZd�0d�1LO��䉇�xd���ϗLD(	6�.D���GOG$ v�!IG�ΗW9ހ���+D�H�g�Ƽ+�=����p��`�g(D�Ty ԃ^�2�y�C�2$9d�{�'%�$(�O�I �iόcR ��G#H�XH�$"O�l�QHO�nq&�*�L��+�B@�2"O44C�n,��,:���� S"OƱ�i�2!i�p�!b��u�ݓ��H8���ҷ{�<`p�]��i��+D��P�B97��Ia4�[
��9����Vh<Qn	���%�4a��~����R�<��I��<T��		��YB�f�<A����.�X��o߇s�L���_�<yV.R�s��H�3� #P�@��o�<�Uc<1�J�g�U�+��U����Q�<���>S@@�C|��a(�HDy�<��$�9,�Ĝ9uHT0톅���@�<���%dM�5�ߨi9l}��WQ�'.a�& >K1���r�ѣE�֜r��׳�yBKʲ�� �"�R*��p�kS$�yK@�����N� w���AQ��y"�y�`�t��h{6�HVˁ>�M���sӶ�d�'E������5?���x���A>�١��3n~����KE*E�X(pG6D���e/�;G�l�U��o�FTH��8D���*�3q.R����7b9NQB��3D���ǧšp���t2�Yr�.D�8��o��©���7>�޹ۇ*+D�D{�Q!x�d.��"�^]�Հ,D���4�L0?hX ���0CR]�Q�)D����,��\iț,�:)A,'D����� C[4XNZ/z?�u�S�8D����
Cn�C�֠E���H�-5D�� � �q��C5�3�LW8G��m�"O��2vp���Đ�\�L�"O�(�7�ڳFm���p��$��aئ"O
Up��A�
�����
"t�r"O����m�oj�U��� W�d��"Or�S��G���}{��K��9"�"O���Q	�8Car���f�:l`b"OuȅJ��X��Q�S��%��q0P"OP��5�^��Rp�	tY�%"OL���Ǫy��59@뇛kr���"ON���|q�עb
ny�5"O(�,�v�tu��Ѓ d�h�"O��i�e�� ��e�8O�	�"O�A4��b�I�p��F��(��"O�,P�Pneba�#�G�-�"O�]�#Í&�D�q����Y�p"Ov����	�L�Ƌ��yctT�"O8M�K
"V]���Y�CLT<�S"O t�B��'\v��EKJ�����"O��xх^*�B���	Ŷ��)2�"Ox��D��/�p����U��4�2"O���C��7��p{�岈:"O��&ɟQb�"�ϛO�1R�"OƸkE��&�04�voZea�<�'"O�ԑʗsՌ�q�Q�/�ֽ��"O�I�cf_�X�2m#!���f0�5"O�5�7%N!p����߉30L �2"O�5kAJ�8
��lX��D�TJν;�"O�z!��$�@�Z"z.�� �"O��A�K�D}6�a���(�
�§"Orp�mH�S-��j�Z��ba"O6T�p�0d����
�]dr���"O��Pu��)?�8BgF�u ����"O�m�˂�<�����$¦��"O�ś� �XXf�[BMW[��X�6"O�@�qȯVb.<ZW���g��"O��@=M�X�*�n׵R]`k5"O�l"��5�ZR֬��Eo��S�"O:\@�.ܓ4{F�Q���5
�"O.|) �Z�yXHWK^z<�F"O"a�����;Z,IH��yjt���"O\�F �(P��4r3�T�\R΀��"Oh�c�˩4���B%$.LU��;�"O�} P̂�A#�����H�C=�t;"O2�+�@M�0��|;b@�tIL��"Of�cA�Z)��W��3$F�H2e"Ol�
��Ja��u+6��.cAjI�""Od,ij�)j艣��"b-��p"OP!*sŕ7\``M�r�&{#��c"Of�`��	R+�4ꑫH�I�-&"O���+-��!�vhЌ\��A�'�<�c�
ÛE��	���۶�+�'��dzD"� ��T`��K,e~@,:
�'p4��B�U3��0@��4Q���J	�'{
ٸum�%�Ԥ�A���D7��9�'(�!d.مr5�0+D�-Ϟ�c�'}��h�G�;Ds�T�AȪQ�!��'���ˡ(�^�L�c˕ΐ�X�'��u�S��1'f`ӂF��*�j�'�J!��#�ƹ�.>*�����'�N�Y����9gL��0$�)�&,��'�����l3-Y��$A��p�(�'X�S'��#p@h5g�*q���'��0�����:�\eXCI����hp��� ��X���9a�v��b()�j��d"O��0m��d��D�`�ݠp�n��%"O4���m��(��R�����C"O��`mF�e6ر�p�n��Y�"O.D C��e�~��U�'M�B�"O���i�+�&���I�!"O�d��Fϑ=���F"�9 FhY�f"Oz�a�k�2<=56�?B��T�&"O�����<wk8[7��)R�a#"O�I'ȋ�g�Z�a����>���"O\]�B�|s�8q�!K.���"O���椕�4�E�s���m5B���"O �0&X�n1XQB�7J0�7"OB]��$<>��UCT+�{*�0"�"On�0�jٛ2Gf=��)��P�f��"O�%�	�Mn�8�B�+@v��2"O�9��3x��=+��"A!ZE�2"O6="QN����`-^A��"O��{���4R�e��"�*W�D��"Ob�;�"Sv��`!�l��@0S"O4��p�Խ�鳔� B���"OVMa5������G�u�&�S"O���a�(��H� +ǬZ��{F"OHxmC�_�|8�#��7l���3"O�(�`E�D��MZaI�QV�q��"O�#w�R�+��p*�e� 4U�Y��"O��!���3n�)ʭK�1H�"OF]����E�^U��+2e��4�F"O��3⫊�,	�HT���x i��"O��Js!�*F�pEϋ�`���A�"O
��Go� t4�iJ���jHTd"OTAH�GX
v�`�/��f�$�Ѡ"Ǒ��<s<��ȕ�Ȼ8}�� �"O����X",�"	���*^H��y�"O�ay�H��:�d������ ��@"O�`��n��2lL��bp"O�(���[�c�P�c�S�5���"O�U�5L��4�na�	{��4�u"O���A�ڭ.�f�����\%�L!S"OX2��S�SN��1��	Ru�A"O8�K���W�4�� �#���`c"O~�Ɂ�̙y':��5J�L� ��"O�eR2�п����Q��iВuj$"O�yA�	?��@����u� <��"O�L�-�
����iV3;��}��"O
9t��^��	(��[�|����"Oh�R�\�p���B�*1�����"O�E�T-����f=۰"O8�B�&��[����{j̑r"O�@)��oF�b�/Ť.JUZ�"O�,z�,OTI��&,>Y��ɕ"O�Đ��Θ���%FL$�
��%"O.d�%.�<���c3�.��$"O�#�	")q	q���?&�ܹ'"O>,rӀ_�h����R�
�2T"O�s"�������3�N���"O�	���:��m��W�5�xՓ�"O�@W�$(�њ�˝k�B4`"O�5��)+@(����{T0�w"OP�C-� =�^��3�I%\N�;"O*=zĤ@�F@P����� RR1�u"O��cA��7|Tr�6���P5"O@��$
�|?��"#@3� ���"O����� BH�aO�?T���"O� ��s,��z�nA�ϔ��	X"O��z)F�9�H�Z��M��"Oi@q�
=��hP�"t��-��"Oā!��Nk�Qs� 4Z���3"O�aK��&@��P�҄/cz5��"OL���,�p��^6�4sw"O֘	�ϤX*=���;>6R,x"OR�����ʐ���L�B0��"O�!qv��oS�\�W�+P��$ʧ"O�� �"�"�����51�����"Or�CKأRL�ĺSlkƚ�(%"O��o�:%�x8��D3z��u v"O����H=v�襂C#���r"OLXQ�L�?#t4�sb�-x(��""Or���$��B�L9�U��"OF��0�G9}XV��O�u����"O�\��܌ʤ���  Gp�=�w"OX9��	>�B�C�#L@k�l�S"O2��1�B�\uR�*Q��NWd�"O�`P���5������	-0ڝ��"O�$;e+R�fkj��cU
m�xՊ!"O��JrG�ˮ�@�0
���"O�y�6�V�Q�A˟x�T!3%"O�B�@��]��jY�n���"O�$�%nI1���h�e�NA��"Ox83���y�(�E�}ֺ|�R"O�D�p�Ź*^�\��a3^
5�"O��J��ڴl�:���N��[z�iq@"Ol�{�"X A�]h���M�n8�"O�Ab䐟wc�Y����B��t� "O�8�Fb
�]>�E&G�l`�\ɴ"OTqIêJ������T�{Gz��"Of�1���-t����FB�b*\z"O�	�`�^�D��U@�!� -�)�c"O�e�G�+/�"���J0e@l��"O8��u�R@��cꏚK��}�"Od�� nE3��s��¶	)RqQt"O��2��͙B�\�B�%�m@"O�<1�!ϊe�lHP��4��"O��P0���10�]��FJcה�(�"O6�Q禌$J
2P�Fé"��ee"O�mʰ���dT$P�"h8-CL�y"Oڕ�%�*x��M���!yJlY�&"O|(�f� �3b|s���D�~�)�"O����C��W��)8�"��8�"O��[�E�ELx��@v*$I#"OVā2�΅@rְp�E$k�D�ˁ"O�=�7�
P�3�]%�0�á"O
��@��d�^��A/�!Jq��Cv*O��@�M�.J<a2��`�����':L�(6��w暐;҉�-g��HR�'��x��V���#�F�W�^��'J���ۺ{b@��L��hD���'�"]k�-�|ȸ� m\�&����'<�X@&�]���¦��nwyj
�'� $K3H�B��P(W팻5,@�C�'&�p9�j$>g�(���0L��C�'��s����Q�C�K�O���	�'�`e#�I�)X*<��ZY`
�',
�yց����q3ܐ(�
�'p�ܒ�Z�0��8Ԋ:�*0��'�x�sA �?1����`����:D�h��9U���qD
$�pd8D�0���jK�
�M(4�$��+7D�� ֈ�b�:^s����D�F�)��"O�xk$I2%�>�S�E�1�Ρ�"O"�� ���P�D��`��y"O�Z���).K@P�"�+��{�"OL1����v=v(��8��T{"Or�Jrl�ǜ V�᳔"O� ��I�0X���V�R-2�'m1OL��֏ܲ�~l����W�i� "O��bd�!�����\A�~�4"O<i��nO�"#,�r���-�miC"O�L ��C�
0�S�b̶W	8�"Ob��e��}��eєO˃b��q�"OLQ�Ϝ9Z <jp�ȗT&P7"Ol�"N�I����Ŏ�,f"H=B�"O�aQ�����(E�¼y6@�6"O��D�L�;�f� i[5?�$i�"O�Q�ԫУ7kd�� "�w��d"Oɚ0�փَH[���2r��5�"OhP�ӑ|.rA��O�(,L�6"O����M=�(M�%IH�(���1T"Oi�!刕>l��+��DKd"O,E�ER��%qTgU�i���"OJ�)�.V�?TU��E.��1;�"OT)���  x1D��Y��Z�"OV�Qc��������!y(�0"O<���$i�4*�`����"O�Q
pLׯ.�<="�F�:S�H�'"OP��G��	C$ձ��\�=M@��"O�@�$KM8u��A!�l�O4��5"O~�:��V�&����Ꞵ^��7"O, �3�ь#��q���N PD��"O�%�q�R�|�HJ�`�����"O���1�

`����P�����"O�9�)��0m0) ���u�!0�"O�H
1��"(  P��>��ZQ"O�Ԁ���~�p��a�� s-�,�3"Oz)��&,gȥ����.\"
i��"O�58�A�}�Lc�A��sRB�	(i�P��¡�&h|��1"	P
�zB��%s�J���D>.N���w	L�Pq�B�B���u���$�밨�'4��B�36�����$���!����B䉋 ��M���*=B*Ya^>�(8�"O��ca��=:�xY�h�3$(Y�R"O�h�3��`"����ڂb��pk�"O�APbR�(�ɴ�}�d�� "OJ�Pf�8b�.U!ӏA2�0P"e"O����{9��	P�ҿ����"O�I��e��A�W)"���"O� C6��)F%�<Ґm�� �}X�"O�*W�$7l��Ӎ/�"	"O�@���o-s̜3h$ƈ"O �#�ؒ{��@�Ũ��Ԡ""O��pu��@U�Ԋ&�4P]BW"O`#BҞ1�|�ɓd�#�>ei�"Ov�6EN;w�|�9�³h���Jv"O� �,y&,��	61�����`�<р [�� �[R�.6?�ɂ��s�<�$��$UrTy#P0m��1d
EI�<�We�x!��L"w�B�Pa�F�<� 䀎�ʡ`!�_bnz���Lj�<����5n �	1%>Ŕ�2�j��<�a���1G�o�Vēqf�F�<i��
%���a�ʐ;%��K���F�<� �Q�6c¾}��MR&�$�i"O����þY<�`��۩���"O����
����UAz	r"O��wE|�`�`TMH�?#j��p"O�P2Eq�P��櫃+>���"O�	�C��E&�L�W�B!^q#W"OqY֢#턘����R�z�"Ol�sv"p���((�5�lږ"Ö�e�6=�"u����),����"O޹i�����F��Fv2��"OJ)Y�&ъ:�m��?Sk*���"OPɳ7# ��X�j�&|��T"OL8�W�+~f �ns�
iX�"OjY�K5i����o�p�$U��"Oҭ�#�� $��!�i��S�l�Q"O䨫2_�|�ji���M�
b\�q"O���eiͲ��i�B��xF�ٚ"OH��(�R���X��ËT2�E��"O3��0���+�EOv'�ܛ�"O~xee�9=ҽr�	.ց��"O��*B�K,|���rA�8��q0"O�`�&�4f����E��\�4"O��÷���!�� E� V<4C�"OP`�Q���"���`�&��O�6��"O"����-2W�Q���9=�漩&"Ob����R�U�r�h1f(���"O�p؃�F�i��er�&�y$��"O�}��#T��J$&��y�F"O�E��Ó{�֨���V|Z8ks"O~�IҬ����7�
5��  �"OTh�%�O�Hڤ\)��\:{F�;3"O���<�h!�Y�S������"D�@�@E��.�8�,H��ĥ D� ��OUI��XQD��/C�̴Q�?D��l��F��&C˛2?��U2D���l[E��9����J*�8�5�"D�� E�3D�H1��U.�Є)Si!D�Б3L�,
q�ҭRb��"v�;D�i���=FG���Q�Y`�E�p�9D��0�ӃX?��hB�":I�4Sc"2D��;��N/R2$q㨌-NԦH���/D� 2���f�`�d�J>DUr$"�e8D��h��Ҡnt�"c,U8h��An0D��A�HVN�x ��.�l�*��/D���A	��i�I:�ꏰ*8��0E#D�P��L�	G㰔Ӧ��Jt&�A�� D��x ��,a��{�F��a�����$#D��+d�P�e�tP�eǗ�%
ܑ���"D���R�E���K���5	e�A�En!D���eC��YX.A
��}UrE���3D��q�+�=-xhp����h�Y�`�2D��HCE��|N$��k�Lƶ�)�+1D���W�K�y�&!H�4�`l��H/D�l�$��5�H�s�䅡N�*�P­7D� ���.n��p�Q�O�<*�(ah#D�X�G%��~_(`w*�3x�Щj (#D��@��V�t�g�������6D��{W��)��H�,�?r��$�T�&D����;Q ����?1 p���!D��
�gӼz��E���\`A� D�\�T���	>+w\��g
�0�B�	L�FL��>
��
T��7(C�	,9��=S�!އ <��A�tfB䉫#2  E�ۏ�h�@䇔p�dB�)� �IY n��bd�l���/<�I�"OnQ�iV ?m&�Ѱh�.44�*�"O���w��Z�Z���[�0^ʀ"O�p"
3�n�Q�'[�_df�
C"O�Cp`K��"S��'e�ijt"Ot�f�Ź.�0T�]"�0��B���y�mIP�����HF�z�JQs2D�$�y���'?��D�W��!@P�2BÌ�yb! 0CP$ذOC2fÖ��a�	1�y�n�gP hC�^Z2���pd��y�šI������J�I�Z�k%�����?��'/�1���L̩�Co߸>�D��'�<�HAHA�B]�$��
ʯ2�Н��'���2�B]���3��|b�a
�'������R��J5����U�<�Sj�_�� PD��
�c2�N�<���}���)�&��)D%s�a�^�<1	�옊F��>9`2�R��Y�<��EgN�y� �H6��� �W�<��:='�i���'\�=�m�N�<Te$4H^�s7��="�sRMH�<at��V����$e�8r�B1S��o�<� �5�~�đ�@�4�0�GA�<)�a_>��v��TᐉQ@�<�t���e1��+��#H�*X�%@z�<A��Fz��dL�9���#D�v�<W�ʀY~`��?W���Hu�<q2ѕc��	`f�=6p���D�W�<a�8'�]2f Y6@���{���M�<�C,I
3����߻&߆p+GK�F�<I��/������J�Z��4����f�<q���1�x��`�Y�'ӆ��f(Zh�<ɓ�D��ԫ�(_�[��p�h�<ae��#.B8�%Y1TJ~�jS�Eg�<��*�s���`O�Q�8��[c�<��5oٶAs�rXl� [^�<�WDR8K��Q��!����(�X�<��(Κ���pi�B��wl�<��Z=4�Ȣ��]�[����Ul�<�@g+�D�S�j�F�\��t��o�<i0 ,s�BQ�CK��#����fXh�<��E�'u�ȰFm<���Kբ^b�<9h�|z�$�@�١H�1sgb�<q4)kײTFE����ِ� �y�<�D���*wĚp�^kv�<�mƌ1VԬj�ԡ���@� Fg�<a1�V�
����:�p��5śY�<a���@����@����N�<iv�\�+�|��]�|3��03�@�<1JZ!rI�	� kr�!Fl_{�<��
Y5,�T������V�8���u�<a��G�?ql������~v0��g�Do�<ѲeU�G��D����x|��[k�<I��a����po؝e��)�|�<�!�ݒ.�D���Zu�� ao�<1�i �j2v)�B�}�Pi@ǃ�U�<!1��!h
��`�A9��	�@Xh�<�3��<��E	r`�tR���c�O�<�G�!:P�T]�H����H�<p%��~�h\���T3x-��ٴo^�<y�K5~f�U��`����Հo�<��	g
T ��c�(df��0©�U�<񦨟m�<�����!?�ȑh�HJR�<�o�>s�8����kΎ�ӆLX�<� �ñ���q� �1�O��Y�=ra"O�I��f�O�D�9!�ȸA�f	�"O���-6mc�)��\7nϰl�e"O�P�R��F��6�ڣ{�*m3f"O���7g��Ԭ����e�
�'�XJ塐0�8Av* ��=��'8�1%��Wn8�y�
�'NL���'�T)�t#ؚRވ�(��M��'@��d0UV��Ѧ��_^p
�'a�4ab�O�ly�@Ȧ(ȭ�Va�ȓ[N��$^�q�F%h %L��=�ȓ&8���6�_�rH�0���!H��ن�O��8�H�(�}��KM(LY�ȓ�~� �J��?��LH��ԿH�@L��J�l�w.�:w{x�	W�
Jv(�ȓ(!��k4(ˇt,��	��@�&L��A䐴��-�3oJ
����>!d��fg^\��g�6*|�ᢥ�_�61��ȓ)�Z#�H�ef��b�.�<#�ɇȓ@�>���S@�
pB�m�����	Z�'����UaP�������=%�l	*�'�jx�_��q���B�n��)�+[G�<A��(��� �t*�W��F�<��9+NX�c���{��!%�<��J�e����bj]�I�����x�<q&����p�ܐo*��m�<��F"p�^�t�D�c�̨��l�<��*Plh	��q&9P�-�g�<���K YgT쓲�ܒ�*�m\]�<�@�W��B��(8ȕ���W�<��,Ӷih���O�t��M3%�W�<���H�=AV�2Gl��9�P`Zю�Q�<!����T=��Ƌ$��="CD\Q�<	V͉vL��&���\�V�a
�A�<A��::4|4��A�842�Ui�<�g��}kR塦I�0����`�N�<����b��\�q��F�����s�<�j��a��,��cA�buJ��@��m�<yvf��o� i6A���Y� ��i�<CeWGl�u�M8n񢠡qg�<Id�#Ab]��ˇ�`�q!���yj%��p	q��*-0|h����y��;yv	r�J�:!16dゃ��y� ~}:Lx�(
�C��\�"���y��T�gM�8���'P���Z��D�yr� >/�� ۡ��E)��ӕ�Y��yr/��d��1�ʓ+.���@e�\(�y���%<Є��ߤO�z!)E��9�y�DU'kn�t�ͬG7�
U�S+�y"�_�Ka�ax&��U�����'C�y�b+L�&�Y���>F_p8B��y�iH���,XT�ĸ<�fm0��y2�I;Z��"��5��Y
B���yRY>t�.�óGQ:3�@u��=�yR�-<�K��$���AHJ��yRd�����5�� n�R�'��y�a��OFT�'Ό�=�Z4R�ک�y��6@Q`�S�b��9����G-_��y��[!I\2�A���)ˈmA���y��G=�\0�É��J`��A���y��>X���"a��yz��!�y���p�D���	�f'�IRB����y"�V��U���M�^m�ˑ�`/D�x��*�WAt�r�T�l��/=D�� ��R֬X�F��|jC��-g�,٣�*O<��S�.|�ȤI��F�L�@���'�$�Gg�:C�jQҨJ-	f�s�'�8t
dk�[ې���@J��C�'�Z$R�� ���Zt�U1~�����'jl��U��� ��oحr6޴�'ŘXA�ǉ�A���H��c06p�'�Q�
&��i	u�A�HD��ȓ:����4�����5���Y�A�H�ȓdӰ}#Q�l����7�^�r�⍄�����Ph!��aFZЇȓJ�4�s��ӃD�T���W�R�Q�ȓj9���qcХpDL�a��'�ؙ��Y�n��Ro��κt/ʧsRY��Q�n��ՅՍqFL�е��PS��ȓ.�p� @D�L���+�"ǣc����ȓ
wp Ib�B2>Ɍ�� ㈟=���ȓ3hqb4*�n=<�d��a����-a�+B�ި[�P� �L��/�`��|�XT���������g��(dY�ȓ4$ɺ���T��u�Ξ+Z���r|�X�@�L�z��b���wv���ȓ_��iZ2I�%ME܅�F(X�[
Rч�#�b�
S �_��R��
�$���ȓ@��;���"*F�9� V- t �ȓ|1P��uD@��%�7�^\�ȓCKL�H�H	J@.�"k��rE��5pZ쫑!L�4�pX3W� T����ȓSl�&cV-�V�����;3Є!�ȓ�`a�d�3
�=IրZy�X���>��q���&v�Z�3&\�d�ȓP�(�!ѣ�46ތ0R�n�q ��
�l���`�M��uh!�WH���_pbY�/�e�V 
Ѯ�5�:�'X�<b��H1V~&,����a�p�
�'����Aa���Fe�3�2W0�|	
�'ˎ 9l�+��-��1Rp�1	�'S�m�/XF�@y&��w@�	�'hR�!�+�� �u/��t�(L�	�'�B9�� V��)j�b�&W��A	�'�xU(����2T"�jǩK��i

�'T|C�jG�o�أ慙DX��h�'��j&/���(+�H�5�f�q
�'�̥���ӡ=��9��4Q��3	�'�a���OH��h���+����'FYbB�5�x�#LʵW�x�'
�B$�dH�p�n�|S����'i\r�3<���	�yp,D��'�V�)t�$?�dԁ�kI*v#��!�'����aT9Ӛ���,�a�`l�	�'� Y�"�͈x�8 �6���^��A�'g� �K]�:%`ٶ���PI����'p��!%Q Yިҡ ���'C���hK3&�]jr�Q� ����
�'��b�7Y�$�c�C(2�L��"OP5���@z0U;�gȃ*�(��"O�)X�!�(��Q�p&��p���8�"Ord#�J�#.�*�a��8:MyB"O~`)BaO�1�����1z�P�"O`)y����QG�&�N��!"O>�9#
�H>5�B�q��D�W"O�����6�T���Z�8�#"O���P��x&V�����F�^}�v"O �ߩ[~���l)@�ܴ��"O� �IB�I�v)� L]��L���"OrM��͌�pY�pI�Lk�|�""O���H+]�H�Ňɮg�c4"OF�KK0�z���E�!q��"OX=W	^�k̎q{��XP��H�"Oh�0��.#v�� #5l:��'"Od��gJ_�@���a�>U2��"Oz�(��	j]��#�{ ^	�%"O�l�$�E�d�5nK�A��Ȇ"O<k��0?��+��BD@��"OT�ZZ�|�K�6,��ң"O0�H�A��	��e/֏�ٷ"O��!��.n�PL��i�b���"O�|���L4%	̝K��I�}&D�"Ox�b�%N:wt�!�a�+P���"O�̒�N�פT�pjO�*��i�"O��T�͌7.`pv��$�G"O¬Q#͘�b�U;�N<t��qr"O �� F�
k9��)��ľ\X]��"Ov��ǅ��F0���h�;B�r�"O�Ӈ�ȭl�zaP�f�9��QCa"OR�����E��]����c�`M�!"O�֛}l��5�ĸ!�"%��"OV����Y�FL�C��޹zН�'"O � !֥�8M� �ٜJs�%�"O!㢎	�`t�d�46���0g"O����<6Β����F�Ó�7D��p���!!�f�U(��U��	ze+6D��R�� ����Ńp�HM� �2D��II��/���rC/)8n���0D�\25J+5���%E� �D(�6�.D�$���t��D��H^�Y^��y#+D��i@�v�*�x���G���z�*D�X��R��,�ŅۂuN~��(D���u�\�3�^UhF�[;
$
�C��3D���ᢆ���iSR�Z�Cĸ���a0D����&�3$f�i׮�>;�Z��c-D���`C�[ ����'�~*�Mp��)D� #ĩ>#
|�䔏,�����!D�l�%#F�S�����a��5P����N2D��!(�-	�f���$��|�2 ���"D�4�Eoƺ�n0�d�� ��ӴH D�� �6*�B�H�2�A`��9D�9bǗ�"��fɫ46��L+D�<z5���X�b��LG�"^2�TJ+D�P�qֵH"�Q�#��&!��=D�p��+��,���٣���x	 1� �;D�,��
�M)�-��5[[ �s�7D��$Lʹ�"Y����7L��{AA5D��Bf�%c �sҌ2 �:#�6D��� �\���0��ђ|\��� � D�dC�$Dx9qv�>P�$+5O=D�\��
?�L�He�m(x��m-D��*�
��tu&X�wAŨ&�xQ�-D�<)�ޠ#Gf4x2��-Z�( e*D����R�{tx����U�h,چ,'D��h��Q��`Xs��:i���a&D�xQG�5K��I�	�Y	FeJ5�%D���T���Q��͉'�1��/D���ێ�T=��
�(���)�� D�,�e��3{��g
J4/|U*�3D�Ȩc� n�t�hQIH�o�TE2'I<D�c��V5/>�QD��~>0V(D��+���9���C���<[`,�0��'D�� ,
�	ҋG���]�[.��"O�<
�Ir-�8���2}-�a�"O�3����u?ڵ;p-�)�)�P"O��1��+u�L����l}���G"O��q�$� 4���ǇL`d{#"O��v�����YQIMG<b�Y"O�	#P�}i,i�I� ;�4�"OB�X��mA�� !BY�`J~�)�"O-I�,�?.���f
R:�P"O>�i���,n����Ԅ4N�(��"O6��3�Ӄ|�DH����{Ӡ��b"Oz�CᘽS�������`� "O:%�Q�ܜj"z亡�_/aܞL3g"O�-���*rn%�@IN&Agv�2"OYa�V�A���BuBЯP��Y�"OF)vFL�{+��f�� !���{�"O�e@�S�tQSJ���h"O��q6�E�Yr��Ɍp��D�"O�|ȅh�T�(2�&�����"O$�@�� �$m(��57o��2"O��17*�	�j��&ˌ'`���D"O��t���1��lH�@��M!�"O4��Mۖ'��%�Iɳv��&"O$Ij�f�)A���AS������"O����ݲJ~�VA�c���#�"O�J3oE Knl�U� -����"Ob9��n�a�x�c���_u%�v"O�Y�q,G�{d��F��|.��"OBp(��F7K�́�f�8i���Ȅ"O����m@CJ4Q`��*�q�"O@���`]�AuJ����Ⱥ���0"O�J���&�2}�V�����qt"O40 ��P�"P��)!���4���%"O�<�s��D���񌛃>���s"O�9R���Ҕ2`E߸R)��x�"OPc�,C?c!��8���!j�w"OpP{*̷Y������B�[U���q"O&����uQ��)3o9����"O1��LБ�X8�u�ڒR=�i�"OR8��!�	`��o��_ ��P"Ot���f_�,���`�طP��ܚ�"O�e��Y\L��
C��]b�"O���&Nڎag�qc�nH@9Q�"Ozu�2$ʱ_U@P���@`����"O"9A-Y�oV�y�f�$5�]�W"O�� ��#W�L�V/�B�&"O>��OC��t��Db�D�%#e"O:��F�0��Ih���#{$�"O&D35��9,H1�,Vj��5"O�!���n�PX��{P$�S"O �*'�dH��f�{J0B�"O`UIckE.`�R �DH�&�=9�"O�+�JE�zc֬
�E�!1��"O8��6�u�PSeX���@�"O�(3�r��3�dΪD�ى�"O"Ex�)!A����LR/9-"��"O�!�F�'<��eM��1&��d"O�a"B�
L�Н���
$-�6�4"O��IS!n�v,�)ת�D E"O��aBV�7����զڕ�R"OP�`�غZ��(���.���!�"O\��kѐ#��8K'���Vm	�"On� ����iyGn�fn��`"O��z��]�	�FQ�V��ljF)U"O� $��V�{`P(�ǻ~�C�"Ojx��˜Z|��F	�(����"O�����!Wg
m�%h�2�@��&"O�9�E��Y���6F�K�,��0"O�%�ØaYb zPg�X��mY"O�S	���.�8�&�#!����5"O����*sA�$*���zVd��"OP����t1��P�c�69�z��6"O8u����
׸\2�C2_��%��"O:�0���;A�|��O1 �I��"Oڬ�Չ^3A�đ!6(Ճk�@�z#"O�!q�B��
�.��2-��<hH�"OB	��J���29�H?r�(��"O�-$��yK��b��=��d{��'�ў"~
_�Wj
`��`[�%��U ��ͫ�yb �u�6o�)ph���$"�0�!�K�q��!U��,}�~������!���.�f���K"&��x`a��+!���5�����	�I�*��ek�;!��	���2En�O7\��2C�!�L��9��mݢk j���+͏/�!�6]��!vOa&�Y���!�$	wI؈�ǟZ|�x2��K5H�!��k�41CVF�jh2������e�!��=j�6��0FX�%87�&0!�$��<,<����:nH��H�)�!��,/�* {7��fH��r�ؒ�!���'3pB���޶{X
E¤��F\!��Z�0�p�=�`����&�!�DZ�tn&�8��FN*X�kA�;v�!�ċ�R{��sL�=G#���f��J!�d�>��Z���%"���AO�T-!��ݞI62PpbaM�a�����G-$!򄉀J���{�V�o��D!t���:!�DH��d�`TJ�1jl>}@AL�/v�!򤒁V���[WlJ���mY0���B�!�Z�)t�2�$�A�dDL�<�!�D�;�P���d̳8W$)@���w�!�D��j�h����R�_;���,K�!�D
;�*�r��M�XhDM�Y�!�䋼&�8��g??`�3�^�>�!�D׼l5�����t�xɊ��K�0�!��ڣ6��H�$�L�@�u2#�a�!��-��I�MǷ������<*�!�$ϟz76��T��!��jeb=�!�dL�`�@�b�Z��G�d�!�d1�>�Hԍ���
�Z`���,�!�$�� �Šŭ�2���3R` �!�D� Ô$��]
fz
��l�w[!�D�Xf�H�F�)	j��@7��!.\!�d��ReظXĆ%lS
���C<HN!�$Y?&�\s�	,r?t�tmѸ?!�d�e�~!��P%$SWl�<b0!�Ā VV} �/��mt1l��l!�dS�A�X�����Xm(�'Kͩr�!�H1OX�I�&1\�� �i��!��\<�T�q�Ct�� �H%�!�A�� �"��U"��29[r!��A-���"�X1��X���<p!���6ʈm�d�^�"'ȸ��.L	d!�D�4d�R,��À0!�xQJ4(�mH!��H��5)6�D 9�'�4}ܩ�	�'Fx�`�)A��@c')��Y҄��	�' ��A�?jX,h$ֆW�B��� l蹳oɼKm�D�����Л2"O���3�E�~u̡�gD(�����"O�Z���)+�c㟅/� �I"O�$�B'̮7���6BQ �^�b"O�c���6�
L����k�d@'"O�}���D/G�ք"��*4� ���"O��r���V��X�ԍK#�{�"O~4b�/ 5�Rc�&�%�"O�I�VM��V΀�BE�T<�1�"O�Y�KH+6��@��3x���9�"ONi$�������z��љ�"O���!��U��!����^mD�K@"O�86�ʢ7{�pCDN�Di�L!"O
	��R��`�d��˷iC��y�_�N%�ZgW1V�^���S�y��U��8�:� H1a�����	<�y�j�:NN��HZ�ݲu����yBL]2H@��QŊ�t�ť[��y��
_}h|c��E1y��EZ$�>�yr���c�<ث��4j��L[d���y�a��$'@L��\$fS|p�j ��y�Ǔ!oV0DR�n~!����1�y��ߋL_�� c�.5�h�iҮZ��y�R(,V�1KR&R/*1�p�q�I��y�j�u��P1g&G&&ObDaт�?�yr��S���bn׬R4B�8d����y��(~$Y�揶5�L���B�yB-�,*W��8aL*0-�$�ׁ�6�y��_� ��(��Y��dpǯۉ�y2nN�kJP(����H�����y��u��X���R�<��x���?�y"nXʈ��jQ3��	�S��y��X�1kd��a�Sp�'g^��yb䅸H�dIE"���qJ��yraL'?,@ҁ.��H<��1�P��y�Y$t�bك���EØ��a
�
�y2B����Г�֞��yaO�y��|wνA�Ƒ ��b�&+�y�K_TJa�b�Ε��@�.$�y2��>q@ԁ#[�}�R����yr)8z6�k�E������d/ƅ�y�'D�u�z=0⃖ 6�AjT���y� X�BGZ�bR@��f\x����[��y�h�:S\�`fA�`�l�+2����y"kǧ$������5d� ���yb�G6T��x��Q�UǘD�cM�7�y��
�a(�*�)_��P����y�ۃmP�9��*@?P�t5c�e��y��_ �D�4��48�.d
`�y�ՏW�J�r���3���gl1�y�aIi�A��m�'{|�{,�.�y2A�cF�p+b!�!&�Љ��A:�y¦J�"��hIU%4@ʈ���!�1�y�5�F�`fn�	L��3����y�$nq+`��7�ڙ	wi���y"��.��0E �"@�t��C�yB%�"�V���Y�0h�Û+�y�h�tz`�	��!挅����yrʓ�<Cl�.�-�nN�N�D���'>V-�KL9�-C���$��q��'��P�,��"�j����S<f�.�J�'R�@ߞ'd�ɂB<a� �2�'��$��.+5"��Q���R(� ��'�di��Hܼ�j�#}�L���� ��ڤN.]u�Mp�	���Iq&"O�E�@@-�Se?�Rq�"O�4�סZ�N�\-:,�M�y`q"O�d�A�'k<12	�
J)I�"O�0Hj�'1d�-X�"O<�k�ȏ�K�� ck[cb:@Z�"O�m2$��-!����+��8m��B�"O�,@�MTp�!��ሂL3�xr�"O^��SlM�2F
E`��\�
����q"O܅�`�)<J�Qp��/?���3�"O� ��p����XwV`�1"O���nOj(CE�c*$�@v"O��0c���`��r U�4|^�k"O�-j�%�1�D��B�h>��jb"OD�b�C�ny�i��h�i1�a��"OH�H���@c~ـ'-�*��$"O�`Z�����u�L�T ��%"O����	͈��ǭ!����"OJ�:�Ä�:I~8�t�TK��Qd"O�J&�!|�2pRT��3V 0b"O\��S�	^2����UUFZRR"O��i%�J�-�y�Oٿ\0�uRf"Of���)��,�«ֶn.�9�"O is����/B�sA��j�5h�"O��)������A���O�"O��7�F	"4K'�&:���z�"Ox��H?X�Ȝ�G���y`L�16"OQ���O�/ʒ��.^&��C4"O�J���?\��҂�*L2
}Jg"O@cf��C�ɋ��Bh�X�"O��GJS?P�v��j�b��љw"O*�'�8?؞ѱ!oVQ��P"O�Q �$L$IK���/`��BU�,�!򤏝K�~\2�B*�J��j�(�!��$�\�aP��DT:D)��l�!���>(�C/á;�\� ��o!�������$��+t�A���H�o!�
���S(�l�����:��DI���e���<W�!�ψ��yB�E���c6/!Z`��y"�2	n�eЧ�)��A"�_-�y�(�<8t�y#GF\R����1#ڎ�yҥ؀Q={W�,N��q����y�3U��3K@�?�l����y�[1g�dڗ.�:��=����y���:c+�h�d��k|0@'ň�y2�B�<3\5�2f	Q�x�Iq�<�%IƹF4T���E�ܽ��K�w�<��H¢�^���p������w�<����,�x�a�-�}�B�K�O�|�<Y�C�OHxx����V8
 	�v�<���M�8���a��}����g�<��"̚!ԝ�cL�Y��(բ�b�<��H� .��Q6(';�a �.�_�<)e�[&{=b]��ć�xP}z�F�_�<���%��P�%dαu2�E�X�<�Ti$e���2����a��ubA�R�<��m@�{�� z�,G�7����RN�<	A$	�3~$C���e$h�Q2_�<Q%B?������r�li��Y�<I!)^�w��}Paf_
o��)�`�<ᡯą<g ��6��\�4�`*^c�<����5���h�ɗj���Q^�<y�z��9����@��ѻ��C�<� <!��(3�e �a�B{W"O��Ҁ$�M�<Q�C�]�t:NxXv"OT
v�I�YG�E�U��-��A"Ox�qb�o���FgVh��q"O
�x�kV;�m�e?<�B�&"OD�+��Z���b'�ӿ(T֐!4"Oh�۰��!YT�qWA�0V�R�)�"O��Y�!�j`C�O�z�%�r"O �2�]��Y���L���:"O�� S@�w���Bo�l10���"O��Q� d1�L����I� ��"O����L�
r�5؅�B���l�"O����̊TG={c��1|�X�C"ORt9ĂջV�<�����3 {��1�"O�<C'Ά�v٘y�B�*#�<��
O�7-�6�r�Â��$a+t��J�!�d��3���k�a̾m�rL���ջq�ab�O�	�4�A6v��Ӆ��-�,��"O��KC��[����%�G�'��I����3.�L�T�A!_H�l��Xt��B䉭v��	���ף=�عգ�b�Ģ<��T>E����'6x(�`*�!'�P��)�OH�E�f��s/��ظ���I�LD�9Zd�>����<F��'���u�E�T����p͍�?�|�"��B妁F��2	�ؙ��pH�-���V5��ā9���&�ē��'vͣ2���
$��j{��dGu�*@�?%>�KN>��zn,�q���n���a��t���=ѷɍ�_\�q���0h�������f?�۴���g�,����OG��賅�P�� p�cK&L��-��'�f��1g�+L��$z�	=Ib Z���'��>���2	�h�Hи"�����;B��B䉈j��H�#aY�g������9rm�B�	i���shK�x՜0��[4{0C�/[o�`�c��p#B����B�/%�<�g��-7z�1t�Qm�B�	C����G�+N������.H�B�	 Wl�%s������蘒U4���0?ل��;d� ��d���g/<�WB�s�<�"�X(Pb�)���C�i��D�P�H�<�Ƣ�:J�2��[#.�"iP��SN�<!����E���s-b^`w�]L�<Q"	G9?�nd�Sn��ǧ@K�<!�Tq����*�_�*�KU�S�<Y$�.���7gY�*��b�O�<�uH*aC�A�=W��(��-t�<�Df8����qG:q7.M��Yi�<QD�s�,k�jO�L���$m�<�vd�'��(�F�K�|�Y���e�<�֍�c�-�N�E�l�)5�V^�<���G1
upA'V�M->4z� �`�<9��ֲxz	�#��k���ykXQ�<	 ���0Ը��!u�x9$�NH�<����*zP��N�*�\��%�D��E{҄N qj�����5.Ԉ1�	���yBc��f��	p�bAS���1��%���(�S�O��!ꦢ��T�T2�k�% j���'
 �7	��dF<��$d��b=��sJ<��W��@1DXFJf�7�ݔ8�@X��k��:%癶u�,� �+�|�����i��L*w*��#1���H�E$��ȓHQP	K�FCP��գ�==���IFy"A�5辁IW����.8i3����2�S�O鮼�S�$tb�A��H@H5��EQc�']?i{�$��<���H�2�"��"+D�� ��jM6�~�xBM ���W�x��)�� �����!R�x�.�� J,�DC�W.�Q gΔ�H�ň�͇�M�a���X�������H�L�&d��O����杠lfH$��*O�2|.D�O$Dzb��(���A���4�{�׉q�!�DV�� �S�ȥa��ٙ#.��L!���`�-��I].,�͟�L��b��6�S�4ǋ=K$����G6_�بaJ����>�J���Џ�+>��Ӗ!�"�f`��JEO~�:O��)��<���;��-#A��� �:�#��jX���=!��ZȪָ�N�	�cA�8����O��M�
�x3���lķ[r�P�i��`�I�����!�'��S�ahW8��(G Ɖx<�P��H���87mٔ���)�Ɇ�]l��'�|�?y���B4sʍ*�E�:@�����ͩ!�>X9|]�c�R��p�W �6)n�ӂ�)���b��0+I, �����8eޤ��$ȸ��Wv|a��Թt�hj4+кu P�<�ߓ=k��ۢ���p�F��Щ�.2���>��'V�dq���O,��N<�@���^��d���I�t�!��K4*]�
C ��x�����M�铒��3���lc�����&fv^��$N&��9��6D��j�Zc�)*UŞ*��k��O�㟨���?�sA���t���<<QPǂ$D����%֭FW��@ϖ�
��5�&��O"�����S,�:4��X>�tj2I�.Pd��ȓ&�v,
���##(%zc�)lo��'�`���	�0��A�����H)����0�c�XD{�7O��u����/�RՊ�e�	m�֌�ȓi����-As�l��Ř��B���OM��O�-Gz�Oޔ���J��0X\m��Bh����+�I�a��D��AZ,���;����ɣ`X1O��G��O�#�퓰�,SVF�T.�\��"O���ֈx��TuNB�&�T:ѽi�I`X��JF� ��V�2��U�4�:�!� %����Ms`V>]أ��JՒ0R�铱n�"�z��$D�hZ'�?^T�6c'5����H-�h{�b�E�yG���d� ti�3���R�<�+��Uf�y��/�x�u; ��S�<Is��P�$�`��H��#�`�y�<!v�L�Z�V��$ӫV̠ي��Cq�<V%�_���16jSV��ܳs�Je�<)���)L��I e��+dʗX�<ɲ/��@2�����݀1i�X�<A*P�R��ѩV��?WJd	aZV���'�����v�� ~���C�i,�y"�#E϶8I��H6w���$iJ��yRj�Hx��p�D��"$��y"m/�t����7]L$)�D۟��	B���Or����ކa���f��\��	�'1��Ӌ��G���0FZ�
����';�5�'�ھh�$�q���#��ӓ��'�*�ʲ��[��b�T�U�Lc�OR����Rt:�!W�#vԴ�P�h�{wa}�O��_`� �2�JйR˖e�~g!�$��';�����>c��B6�ǹEi�O��=����C׏L��َ"�X�S@"O�8R"G+
�ܜ��E=���W"O*4�F���:�H�w��2��6�'�!�7kH?4�Zh�#�g��"Q�8��I?9�p����|�3cAݠg����$5�I۟`CקIg�^���DY�^�9�w�'D��竘='q|�BR�����A��'O�=� �����D/'A�l��J��G�H(d"O(Yd䜕
)$���I�M���Q"O��Q7�ɓ_�@pr�H@�#����"O8�I�h�f����@F*M�\K�"Ox�$�"�Р�`�Ev���v�C�O��8Z�"'�0�C%�4���X	�'Q\���N��ځ1�/�<��RN��O>�=�����s��IU,j$��i�����*��I�v3���pE�o*�\�\�B vc���MN���Ĉ"cy��L�}S�����aښ>���9���B���>?��\j�de�X Z8.�Q���On�T��C����@
ƪ8�� N\4%�&��ȓK<�Hå�U.Ț���S*m�X�� A�x�!�<�z��#�Ϥ5�2؅�Kj�0`d�F4V�$\$aS��ȓh�4���%�9i��d`���!D��}�ȓ B��G蟹`�L���!M�`��W��MP5/]*#�IX�Y8vE��y0v�:��-��@�2K� ����L��@�D��"�>,h� E�F��ȓ1�y	p잖:`A X�,���dP=Q`n�o��T��oW3g�f��j�t,�KA�k~���/2Z ńȓExe�Ġ�F{J����)��p��t��m`f�C.4���x��̂@�`�ȓ ;2����}F���dE�wЇȓ;Fl�bW	X$v�Lhx@�1�l��ȓ1�V��D`�;6�З�=W��,�ȓI:xH�,��-��K�
�tՆ�|{�q"3d��Y	Pr�t�A�D�y"+^-Z�x�pG��;G��Q��ya���� �EOܜC�̰k�D7�yBƒ� ��Q�#�17�
=3VFO�y`�'Z@sCT ����D���y�d�	#Y�,Х/ٸf>����5�yr�Ī��1OYZX���'dŜ�y�}����;�$�v���y�`��V:\A��M��.�H� �y"��({���:D�=f�(غ6���y�@B�����,I�
8����)�+�yR�Тd��H�ǜ�mjН�R����yr�	
��A	D���d���2Ŕ��y�J6
����N)Y���"e���y�씇=�9@k^Ll���b� �yR$�"d�l�V �3�<��BC���y2�I�o$����a^>7�2�*���y��Q�_>\Р@� � ���ď)��'���q$N��i���

0��y2e���d�u��D�*���(�yR!�./L���c�f�6)2!��-�y���=i,z�{2��m6lt���ڥ�yB�9h�FE�#!š~����Ȑ�y⋞�A.�Bď�o�p F��0�y�Tg�Ѐ�v�H����v����yrGP;c��ȣW*_��N��C���y��ՠNy�+�
 #*e��"�*�y��L�cfp��Ȕ+�6��A�K��yR�^y�q�K�/~ L�Pe�y�	8"�č��H�w<8g�[�y���5� ,����?�<�;�AQ��y�!B�=ߔT�6*��P�IF����yR��>$t��H(6�*�B5�y£U�+�b��W
/��uj�ğ*�y�i��9�H�-$^�S�bS��y
� �<����=L��mX�d�e rTz�"O`��۔h!0\�ŔQ0�ٓ"Oh�v�9���D�]L���$"O68�S��R�|1�I�!g>F,H�"O�2��Vט}��,��3�"Oб u"�uK�|z�n�]�%"O�D8�n�v��2��� ���2"O U�%.A�\H��HGo��P�
�	T"O��j�#Ҽ2Vv	�T�S?2�\T��"O�����:��m;3���G���s�"O��VFU�>H()���Ƌjq(��"O �paC�@5�$����OD��s"O
]���Q'=jYx��)1)�[�"Oxd��n^'Y���f�#jhka"O�4����hOJ��t%\'�� �"O�Y"BmC#��l���D��&"O8��u��.Yf"5QQk�Nd�xk�"O>,�PŁF���j��\S��
�"O@�Q	��%і�1}��3�"O�y)G�E/5������U;t"Om���m���c�6J� AiA"O�i ������KC�*�.��0�iF\л7�'��`����(#���eN	Z�f<�ד9?`E��6?�0�.6V��Te��H�P
iXB�<�	�0n�J5j��̑��<�Q�NX
!؃�(���ˣ*=|�d�3tm�j���"O�Xg�ӜC�j���O��2�)^v�qO����Y��c��н+� 
 ��1M�Ν��,%D��ӌߑ�!�/,R|� �IE�1��1IA.�O\���oP�)����M�A?U��',�]S��PO~�lʋ>B��# ZD�p���1�y�I."�) �O��m��a�dݵ��'Z:	[W���d�Š\Q��P��Yb`V���J1�y�iʨ�MaUdVy��sQ% ��y� ��;���3�J�E�uIQʚ�y���pHj�ST"�:=Z��/�yb�ǽy����A�3=nͲs�K,�y�_tV�%��@<*��8�*��yB�I�(���jBHտ#�t�e �y�U%�*��5���gž�y��@?S��waDS;b�zD���y���>��|3�GK��|J@Lѯ�y���y򰐊D��a� |j�Q>�y��9:
Tt cO��W؈����#�y�ɍ4tlu[F�ŦK�f�kf�\<�y�_��y��-|dx%�N:�y�m 9A��U#�eu!䥛��y�� �j%XTy2̦d��*�(�yR��X7�t唪X( mB�oϹ�yrK�v�X���.�R��LҖ ��y2ep��ӡC©IC�����U#ڰ<)�c�S���Op��`�_�N�" P�+�ި""O ����A7�%����:mFQ`� [2mš]v܄�Ж>E�4�-^/�=z�J�D��d�4�y�iS5[�Th�խ!w��x�P�^�0]���O
�St`����&>c��{�s��԰s_�J��@�@n)�O$�CboE5!倔�p�ddaD��f���h�!QR@��Ɩ��	���z3��O{"�S���7C�鳰��!��၉��=G�e$�[?�q2��z��ɗ2���j���x�� {ƞ��y��,t=B�כ|��	�)���y��G�B���?R��\Fnt�  U:w�U�(���i��m�'Y�]�O��!���#�I�M�E�'��h��o�:'H2i��I�q�V�qs#R�#���q)@3���!�*T2?.�2���|`�+.G�T7>)ؠ֞?�T���8�)ȶ>�:�����|�o�	Xvh��FִP�	)�o�?K��,e��#|Fraáe������Ԯ3S��)�W��7V�) OJ|��h>� ʨ"�j��:HLcF/�73��s�%3���ڲ�B߀��c���@��@j�٨	>��uHM�BU�wAr��؀cS��R��A�s���h��xC��j���'�Z�W�p�H��O]��A�	z��aU���Hx���l���w�:��Q	A���etdj�
�O(�&n���(D�c\����j�ʬ1�.�0I�5)�`={fa�F�Mg��`Y#��e��pW>�SC���oG����C�u��_�%��0 �K�j$�1B�E�J_���	� "a�� H>m!�9k��l�T�
�ݸ�"�0C�8�)p	 �}�X5� ��j*�4M���铚�Ԏ��$���`Ś�p��		�hO�C��I8ol8qƁ�Xv�R�^9�d�֭@�6%�6�t�R����e�v ��Qf�	F%�Ei�~�*�`$��R&]J�%�3n�s�V]k�k�O�m�D���:��h�(��"��
r�ݗI��=�N�~��(T1��Ȼ�Wg���4cG�e?ֹ��L=~z�	I1r�H��'q�Ա��L�h���aO
:]%c��Ϝ9	Ȍ���	����q�Ѱ�ug'�6���b��-��i��q��$	�\$@A�ŋ���3�G(�O���SĎ;��I��l��`T�q&��h�ܹ0���M�X�31FT3l2���n�J~"�L*a7�L�5����d͘8H�s�m�l. �RG��#UQ������@֒}`�&B�)qr��O;��ƃ�s�$,�b Jî��ZV�	".���v̉-��g�{Ra����E� 4�.�P����t8.B�!H�s�,�����⤹G�$y#�0 ҂��,���P��(/������ʂ /a"�el^�At�!1��P�A�cQ&IQ�6O� B���(���diP�y"ȡ;�'��hb�ʑ<D\���·s������'���BI,};�bpJ
�h[*��Z�R����烊 ��Й�%	+�=�<E�t�Mpa��!Y�Z(ܜ��X��On`�Ы˟���JI~�c�C�KN�M{�iX�8�ԍ�N�L�<�잶��
�I��2����cy2h',��&�,��'�1��� 'R<��,BA�3���`Q"Oڜ��	�l�u�JйY�V	1b��(�$��!q���&�"|�B#Ws&���o�d�T�*1��S�<�G�>}�B2e�هe�!BFky���2�{�lV���gܓF	P,2�aW�#���2w�5�����	�D@��/߃VEABC��.�N�q���%Hu�'�>PY�_	�̂1gX�%��Q{��$ݲ}/xؓ놝`O�`rg�a>E�'I�&��iV/P�f�D�A�*P{� �qr�)�O��)SEJ	޶��E(��V�2ygY�p��"GN����ܤp�\��'-�v"t ,��ɞ
D �m�邬��� 1���!��*��)�Cʫj؁�䝓d	Ҹ���^#m>����f�(/J�)���j�	M�SX��2�aލrda��<����Q��4M?�O�B�!HQ́��
Z	G>��R�E�.��	Q�^��:E*:lY�n*�H�D{�&Y�xN�P#bN�(4 u�Oo�'��-a3mH8JͨP����;�B�Ivh�6�R��|�U�~�("��A7�J�{BNWX�q�n@.b�Xr.T�3�!
b�#?d)~b
�kd���$���e�CEڵ��fA�FC��AVb�p��ԷDOJS�[%<f,B�	�*���&��5�h)�FB�C�6�����Ff(�[S ϗae8�H��C��
�f�4�h!�B�2��*� �s@@�Zn2d�@	�8���!9 @�X�!�O��Jtg���dsS�*5!2Ō�@s�, 0�4&�1�/�&Y�T�OB�'�B�0r� ���)J1n�(�ҍQ`[v�H1�VA?��ʰm�& ��ċ#��#`�[}ŉ�2bn��pb����ɘ��0O��!�i����R�1N�
#�-ט5�VC �<-Ic!D�����-e�e	�H���Lքi��ʼ;�A�$&lb\�� /N߄�jaH�F�' > �P�S�O @����W��]з���R�2��( (�����3��=�*�C(e�&�|5��'���O�h �����m�bɓ9��������M� �>�iݹӐ<\(m
��Խ:W����4.h>xT
�Y��C�^���E�ȓ{D|k�"��{�x��ѥ��>)��^�؂�Ȕ��!�Q�B���K��,����^�d�7 ϕ^6ep�g�5swa}��On����I�U�­�G)��']|4� .�)1�8�k�j]���Xj҅G��ְB�N3����-4��!{���<$͘C�Ԇs<����!,�Hޱ�| �%&S/(�Υ�e@�)�$*+�����o*o=�4h�����8V�~�<��'O�DP&X����&�"�d#���LSDu�'��dж���WH UrAhF3p�g6Av�p
�j%T'�	�+��~�'�	U<"���'L�t��DǬ����ÇzZ��P���B�y�I����%5(���2��h;�/y'D\b�d�-݋�"O�,�d��xҨ�ك"�v�=��Lb�DE+���N@d��C�7���C�� ~ ��0U �#�xţ��'n��3�8>af	�"B18�(R�N3� ���FW"*!��K"W�@=S J�9=db�Ϙ'&�ѩ&� 3�D��脻G�x`Óh�9W�R?����|s�� DIr4n�k��}{�D�x*j��u�T�D�q���6%|a|�-3ux���f��>)�ŊW�Ԅ���|P��_���S$���a'l�� �"�ӣ	�*�I፟�\JG_�!C�C�	�#��T��,��|:�ٸp���R�H��ʅ?�>,�w#ZȼM�l`��v̧���$"Ө\�����3D���	�������U0B��;Z��+5 �&�iJ��N��'&B�4`K��ϸ'��0��`lu�X�% ��Qy��k�H�1+�	8��t���$��-ް �@ �U@F����c��B*=����	�8#.����#��SFo��@���ړ���,�А!*O-[�Oz�4j#�����'�����-K��p�wJR�h��J�'����T,�fs��yG��hF��@�M=J��`�g�t�Z���ψc\P�DD��J��nN+]��z��I��l��
��=!��@��&��4��h�������G���y�R�&�R� ��b�٣U�ϫ��'���zg�&�h�;sZ,	��	�'m�uQ�I�R.,C�ɷay>dKTF@��B�@Q�1�,\K6�´AmX!,O����Y�� R1O&da�cؾ^�.)��M T��UEϕfJ�8@K��v��ѡM�ZP�@Q�A�� ��ͅ�	�{I�@�uK|�F!�v?��dW(��ˁnG��?Qb�>u��X��g�U7�4�N�{�<��*����y���4}T�!�À�\��DsX���՘ǈ���r���T��L�bF>QQ4|Q�*Ot�J$��:ʅ���>�!�	�'b�U�W�eb�
d�?ftH��'�~�`w�x �t�3�ſ%܁�'��݀��g>�e�NA�vM��'I��!��-i�T�Y��Z�E)\a��'�`��$�U�_�*��`�8r4{�'��i�NC�|�f%H��²6�R)�
�'�Xi��U�_ظMA�)G57ﾥ!�'T^T	�[���f�+&�Hr�'���Q�/��N^
��q�� �H\9�'��P���H�L��Q�aP�yJ�:�'���ȑ*,���'��+ H�2�'��Ղ�@`�I��HG($a�'�d q�@��7K
C7TyB�h�f�<�L�91��2f�	��h� �T�<��k�<jVE��'���	w.T[�<q �z0P��]� `a�W�<A��,8��Y����0�`�X�<Y�]�C���+��j[^��g��~�<��"2"�Rըg	�:rt���l�<QG�;P�M��lB�b�L���fMm�<�����5Cu�c�4����cEB�<9�jQ�69椊��f�D��I~�<I%�%y��́�G�'8,�5��W�<�ҍ����.O�y�z@�5ƙH�<!���R��@���θb�@D�<�����rچX��dZ$A%|���B�<��`��c��,:wN�V[Hk�N�z�<9��;���B�,Nqn�;��x�<AGپw�P@P��^y����K
L�<����_>21�D9�6�
$�L�<�)��w<:1��*E�T9��
o�N�<I�A�8��I�A����W�<1F�����rD�T��]R�.d�<��lS�?�B@P�ۈ^����4Gd�<1�㖊6\ȼSA�C���5K�g�<AOΖ^�$h�]+x⁩�c�<QB
�2w�إ��5|w>y`��Z�<I��Z	aT��$ڏI�,�H�EWV�<�4�D*5S���̧P�� ��V�<�� �R%�x�%�u��0��^�<Ѥ��5τ�`�хb��0���W�<� ��ӭ�N��y��� t��d
4"O �qs�+H5D�cGJ�?qz<Y�"Oju땉�_ל��X2h��1(R"O��B�� �����_�ZW��"O@5*�!}n�[��R���\Y�"O���7��ۊ���ɾO�X
F"O�Ѯ�X��](D�l�1��@�<�@ˍ;~�Hp�Y�{Zx)��F�<�Ղ\�<px�+Ծ��X�S�C{�<��m�T@�KG��2K���bř{�<�&�ٳgO@X9�L*'%�=:&gLs�<�2*	k�0	(���<ܹS�FD�<9#腓?b��q�_|O�-�CA t�<yP�>s�<K��5RIV��\�<�'��+�2�a�qNt���O�R�<� �ߵA�L�b�"R�̒�V�<�FȢE�ȼ�q��0��Y2�i�t�<A�F�)�������VY
�!���Z�<��P=F�Խ����7}��`2��y�<1sf�/&�<ҡ�U	�(�i�u�<y2�R)�N|ӗ'ɵ^����Uq�<��Cާw�0\v-��qZ������V�<y��J�&`�$��e.�,�t�Td�<�c��pk^U��N���X�bI�<Q!�-k��$p����H��q+}�<�7��EP&�w,C�n����WbGA�<y��A/P�հ�g�=(g8����M|�<�E�.w��ш�D�8LV�9���{�<i�MY�J�[�G��l��d���Y�<�2��F>�����(�2�	�'Q�<�Qe�=��e�7�`^�5���FP�<��HD������ D&� aKR�<a�E)���rN<K��`&�[O�<	Dl�(�U���B�"�h�#�s�<��ϛ�O�T@���<y�=�"�s�<a��%F����D	�9��r��m�<!r�O;�L���皰�L�C�#�m�<�ÏD2
��ˁ@�T8R-�M�<��ĞX�0��Q�)J��XȆG�S�<����`�����@�X>���U@�<q��)<���rV��h������~�<1��3"��Ս�Ae��p�m�y�<�$N^77^�yE&r��8�Q��x�<�� ս/��y���ȡJ���9�p�<�׀��
Y�y+ҩ�**l��a��[�<AB��5=��P��n(8�"�~�<����,]�1�ܦmP!�a��{�<���	we�	ು�@�)R�Vw�<�qG�r�(A�e��U��P�QCK�<1�<���d��,�Ar�WA�<A�U�W�Ν1��Jb8:�CB�<q&DA�*��E�!!��]˵FF~�<�r�G,�r��\H��KX\�<��׼"����ꜜ:d��Ye�Q`�<a�E�0�|�cU��8"!��f�<�V�� ����`T>s2��!'cc�<��`ŕ^	LI��o!�`�fn	`�<aC�H�X���t�۽H � 2��t�<��!ЫuL��v�ߝ[��� A�Y_�<Q�F[�`ȷ	�
���8w��Z�<����!72P�Q���$��e�d�UU?��"�<���'��b\��?��G�\ wEn}�-��~�B� �*�On��EBE�WJ�ֈudV(c��y/�����\l�D2d8
�ׂ(��*Z8�eSu'R��e��⟄S3ҐW�|�ۆ��*!���� 4�`��N�]Wlī�h�zڨ�Y�X�Ao�#z�}���'a��(�	ՍLK��#.G�]ub�@T&Ȍ7�D���� :�vp���O���rhM�c*̡QM� ,ʦ�Qga3 H�sa&B\H<aT@��n����ʏw�q�E`��ǻxc��H�@ۆ�T�J$ 	 n���>��O����%� V�ܓ(��q�����X�l�z�銝^���[����r�(��A��ZŰ�{&�P�)נ ?,��L;}r��9����l�%$Mލ���4|b4�?�Vcώ C��?MB����TK�,%���d&�%�14��'t�p�d��8]�ڈ�剉}��P!�/F�%*g�V�H�ЉXPǊ���d!� q�j�D=�S����cq���g��1�G66t�H�C<[��	[��'Ò!8W�G?a��	1������3��g�z������K����<�H�S�G>g��	�}�v>����,#�l�i@`���{"+6�bl�7#σ[��G�[��U9��ҹT�$!�0�ܾg9�LJC:�<�kei�6��[�#�%5�T����O�����B��Xή]ip��K�Kߑ���Y5) -�b�|�3���d��J�IN����1;`��+.��툥�H�z]�es7$ �M����-\Ο0����6vBaz�#�Npy{5��&/6|��@�����[�c 4u�a+F.�0�mZ�MfQCE�%)9n���ueR��dx����:��6JQ��p?AD��O�J<Cf�_n"�H��$�j՚��J�g��7�Ļ�v�pD/X���?� ��ޭ[��ɍXX�EiY/\(�%W���>��EQ�]��])��%�S7^|@�����ZU�uDU:O�h��Oĩ��I(q��%>c��)�JؒO�>���NӬ~A�bϩ�t��	]�q�r��Л>�}����PȮT���66Ȋ�9���~���@$���J�*`��	�`���j��I�I����	=���'�T�y5E�$&|E�ɚ[
� �c���ē4�@\q�ڙp���rT���O/����>�p�:%�rs0dZ��(m��dz��ʿxA@5'c������e��b�"|jր��jN0M�s'Җo':�J��j�'��D[�Ɋ�:�q��4���+y.-3��3�����"O�0���X�h���&�["C�Ҕ�Z������n��'XN���H�',}�����'S���P#Vy<��ȓy��qH��p��#l�e����'"��ja�؅0�ɧ�ʹ������$uA����a�aJ�"OԼ��F	�-皴8	�7a`Y��{���u�Pr\�ϸ'{����!	�.W��y���"��Ya
�'������:��0󓈌 >�l$����� �S�,�O�գ ��t�Mђ�
�(D�D�	�UWƁ3��)�F� �S�|�A샢F}x��2#�`�T��z����a~$Y6O�n�c�8
}�|��@�Z#剣bH<�y2M^� �b� ¬'�
��"���+(��X(�/��}Ɇ�U僴b���"O�@��"JÊ-0�ˇ�@%��*�"'�05�d��rPj��D(���|툴(��W�Z� A�f,r"��!�2�'m��n=����B�r�ڀ�!t*r���0�"Lb�릟�1��C����7�"Y=xE��I�{�'z�Cec�,9���S�"����$��H�V�̢I�V��pB�_�TћS+Q�]#�qqG�Pd7@�[G���*��V
oY���dֆ/u Q�A�Gp�3
��P��I88�&�%Q��eXe�ׅ*r
Y�a�\Bn�ce�G��ѶQz�Ek�Fب}�L䳄�I��y�+��C����V
�wݔ�p$�a�|�[:i� c��	@N.�8�k矈��vJ�0wݖ�`$dC�y���|Zh0�p��3��yDO�0>�`F��p}����7nx��M�!�ʝK@�l58�"C����t@"�]�f`��6���?��p�!���a���p�T��.u\�$#�eN�<E�Q���O\�v�Y�-sV��J�*О���BIY,�`c�t͂bY93"���G����nV���߁yV�UZ���[�v���^�ȣ�L�"Q@����w����������weU��$�{R`Isg@){���	�'�.x�������siK��d��"T�m������n6E���R�B��W�	�!��'���O���.I�
�F�8�;<^����'HD�f�Őq0v��b^�]�`7�@<!,��+5,�,(H! �6�!򤃧z��p��`��`�a�/g��I".5�a�gBAW��e� 韹2�>�ҕ+۳�Z���TSp\h�V�>D���mF��%��ES����Jب+�t�����Y2<�a���x����qO�܂❼y�����F.q��%�'�����b��X<� xĮIl�b���a���)۵#H�D���jj؞�iC�
FN$-�@ϕ�~��1V�"���e��'����/޽5â\��'j�	>�O2�(�N�F!�DO�����Rz� a���
�	�v\١'BE�0 ��F�k�O�x�s�B�W�^����,���� �!���'��L�u�$k(d]PEG�Z���J�D�� J.��$�D�"�K��8zL��aAC�"dV�G�f��DE��v�-���Y�,���*KQM��I
��L�F i��y�`G\�{U���D.5\��;�DT*zd�	��}� � �mАX��$m͊E!�ߢh*��&��I�D�2\�E���ڔ&1V��s�l�X�mĈ'y!���
M	����
�&��"%ދ2�b�P�a�nA���'�8,ڃ%͂S�y3�B8 ��Ţۓo$
E W�T�Z�R�䆞p��<y爞���TN ��!�$�4-Ԍ�6"�,�U.ٞ�qOp����X��q�F�?�'R.`��B
4M5 &nB�eT��ȓp����T��#!t|�+� A�w�RYK�܎J�$2bW��k�<Ѳ�R� ������.-�ؠ��p�<�FG�*e�h���E�$+>��(f�1ivδf�oR�T���'ed�2fO/#�^�sԨ�,�X�B	ד���K�%�^���4YEd(3s��8g�,���J��܆�!Y5�"�J-��zc��=A>��=!�"\9�H�H� @���U�/m� ���C�;���F"O�y�2j˽J���"�"�"a�K.�����!zy�-�m���-d,I�w*3y�4�a��f�!�W_}�T�&k�xS�<F�	�t�x���G�$n��L�gE�S؞��^	J_,�y&F� y
0��D=lO�@1�����[��=A2f��f�0�r��>ax��ȓ;�Tu��O�0�x��K�R]�?YV	ԪJu����	�}Y��*��T�E��Pӣ�#&*!�_:>��;���x4Q�ݫ~!򄅿4��哵bӮ����EƱW�!�D���D�t���|Hy���*�!�RTx<i�(��U���tƔ/(�!�DM�^lN��G	J��8�'�+U�!�"9���ӏP/i �+煔27(!��T�1����
E��ع��>6e!��Y��(	�&�8�,��"#�%U!�dI(��+��ߝ	��e{�`��V�!�ĳ`8�X�	Lf�hiI����]�!��|k@X�c��*�v�2�-�!�d�<iѴ(#e柝t�BQ�'N�1�!�$��[�IVn܊�x�Η�3h!��-,td��"�۶��TAWlD7M!�$U1t`f�hĭB�O��\��M%:!�D��t�^�[��B�*# h��;>�!�Ą�W�0=�ҬŽ=�Ȑ�G�C�!򤗉c�p����{�*��Ug�&,!���$$Y�do�9e�(��b��7�!�D_�+$L Z�cO&�B����[�!��� �a7��n�aP�p�"O��QC�4t�$
Ů��
`ʷ"O���Q%Me��5FޭP5~�f"O�L32�]<0�ʕ3���/L&e��"O`���b\�R� �r�n�/	3�D"On!���RW��-��q�:��"OJ�yF�F�g�\��2�Y��P`""OT4R��˔b6�6Bƚc��m�""O(`bD�aA�d��N4^�����"O���cՒIZA�P�J���˰�(x��۬<?J	pd�7{�'>�A(r����B�Ic�u����C���*7��a�T>����ێM3���N�(>�,Dx����;�I3z��D�2���heb�1d@�wk.(H�OfD�gKXn~�哢P�^�17A߼eD�QtO�G��7Ͷ��SFaD�����#u�@ם�47�M��D�T����J�p�$L��O.)�)�'�l#���&[7��S��E]��p���ܲ��'?%>O�y:~q���80��r㏏+���Wg�I�W���>��`�*:B[�/��W ���9�MQe��ܱ`�Oa�� D��Iˁ%T`�@T���-k��i�qO�)�S�O���c��aq *Z���3];�c���h�t��g}����"�UK'N0���dh���֮N�bP�{���8<�|ٻ�b�L�8�Q�&D����=;*4�Ɍ{��i��־=z0�	�&�\0(��o���p͛#��I Y��=�)��c�	F��0�(�LԂ5�Y��b	FxJ|�1C��ۧj�D��I �R≪�#<�~�"J��{ L� 	1��c��s}AJ��O�>�qNH�DZ�:�,|�>�g�e���&�i��D���~��D�?��#�G�Kff�ʧ���S��{2b��>c�	�m����D�p>u�*T�Ist���&qb%�<i4푑�@0�ԩ�|��0E\a�%��*�z���S�w=��I�YS������
}1�S�O�\J���DQ��{d�m���� d)rM��L�%~B��S>[ZH�0��$}Z8(V�dSZH� ���}[��C�A�a�t���(E�Ջ%,�	/���O�P��BD}?q���?y���O���?1��LU�mLB́�߁p�L�7-\�o�V�m(9���3 �C	�����(`��fɛ]��)['�D�v���	�K�n�go��a&(��剛J<��t�%q���To�<e��B�I1X������ºT�h���^H	�B䉸>����3+-$�Z�&0Y^lC�	(CBi�#�6[u���fÚ�#�VC�	�S��B
^�����l��?�B�ɦe��YC�kB�t%�q�4EM+��C䉸e��*��ån�R܁``�=iZB��iG
�ѣ�	�ts���y4�C�I.a�QH1�4%
l��#�t�B�I�'|����m�)ږ��Q��C�I
G�`�'�ne	�+ǱK�pC�QH4��� �2%J3M�dPC�I�Vg�`����\�Pq#��)��B䉖>�z0@���
VO�}S@bܱG�2C䉅3�����,��-�����6	6B�	*�f�2ff�N1��(��.�B�I_��ƊD��)�� �B�I���� 3c٦eE�p��EQ�8B��)W]����EB�!����g͑*-2B�	�$S(�����x�x��N��C䉼(�ԀB�I�FV�kW
$5 C�	1=�u+�M_�D�K��Ƹx�B�+>�J���dا��J"�Ǹ&�B��$,�z [(�k��]09P\�XA*D����xG�2��
?�����'D��B�oޠb!�1�/mL��G"D�� 6"�&�H���*նq�&�jR� D�"��ڲgiZp���bm��9�$1D��钇
|�.�JPA�~���cE1D�H7�Vtv��-�"E5� �M0D��z�K":6$�V�_�7���ZD�+D����-ƫ,�>p�n��4�P��=D��$ŉh�f���,Vt��@0��=D�tK��R�M���`�El̔i3�:D�TID�T-r�)ꤤ�rhY��6D���5A[!���q��T�~�P��4D��.��,z\u��4\�ؑ��1D��*����m��V4�A�.D������7td�ن�/�,�A.D��H��Q�k�2��s�@�yiB���?D������&6�t���\��Π8S%1D�\:4��<A��%�P�}d�p(a	.D��B��r����Ę<N��9s�?D��@���>jԌ�#	L�y�9�:D����,t�x4��U��	=D��BW�A�2�r0p��K
vh����8D��kfa}�pۗ��%��ĉ'7D�� � ؑ��L�d��7!J+L7�}C"O6�J����|m�Q�ߊa�`�hT"O*�����=b��2N���B"O`��Q�L=A�X!�L��*t�]��'�A
���n�V9�ek>.�ą�
�'ܮ���/��h.>-�� ��]��'���J��I�*��e�	�.�`%(��-5 �^
Ha���C2QvEB�'h��U?$���`%n@�Y�D��
�'�h�2�P6zt����&�J	6M�
�'�LL��E/��-X�C�P�8��'��{��P�|z4X83gH��p}��'���{pm�5*x�j�`I�X�����'@���6��;uae�HHN��ȉ�'���1�ёx����=B����'��W�o}l�T+��.��!	�'V�lڤ1s��@�
�>�,Da�'H����	ãY��*Aʎ�p���'8�� �Β"`6�Ґ.̑��a�'�p�ш.���Æ�״4��'P�A��V�V@�D��"}����'P�w�^'F�.�!���Y����'�}cEjϦ6k�qI k��L����'��A0s��,ڼ��dB�znR�Z�'��󕈏C;ba���Ĥ\�m

�'�p;v2�Έ�"��<�i
�'Y,�CҬUdV�`�ݭM����	�'�tX��.��y�@�"Y�V4����'�j,�&�B?6���'OK�����'���s� +0舡0nH�H�:�'I�hj'��S������>�(�!�'��X"�
�X���� M�ę�'r��0h�+�I�E�""8���'Oй����4}5�p�i�������'���;Ҭ�9K�J�n����	�'H�]H7�R�8���Qd��u���'d�(��Հ;D�eX�a^�b�:0��'��8�`GM=j\�	×�Py2��	�'PЁڳ/.	���C�C�>�p�'�Ԍ���
HUu��?�0���'���wo�1^�8��
"4�:%1�'C6Y)A% �(�i(���1k<0Y�'}�,�0g��IY
�"4`N�Q%x��'���HD)Ȓ��SE�N���
�'l~q�p�R�<L��f�@�@	�'-|D)�M�L+@9�28kV���'�� y�c
��b�Qa_�X��9(�'�J�٠BIh=쀘��Fh>Z�x�'�*\y�+M%����N�_�D� �'P��������IX�X��$��'}8��tO�9?܎�xF_��\�c�'�}�Q�Q+��8V
��kQ�'ܦـ�P�wX$�P�����p�'���!�H?E��y���H�w��
�'�XY[���*d��9��/jZB	�'��m3�֏W6�D�f�ya�	�
�'�eX��1��ɉ�j �Gg��'�,(��1\�
Q�ȧ@�n��'��K�%Q5��бg��?�Y�'	�և; 3Ј!��ƀ=�)�'����Ç��!��LP�l�^�:�'؆�ےEB�{V���a��d���
�'@@�!�ધjH�(�^���'�V �����'�bm��P*	������ ���Ǝ�0����<���"Oԙat��B�,�:�� 1h��e"O���M��%��t���)�}Ӷ"O���r�[
�<s5d�6z	B�c"O�<á���)P <��E��Z�i�"O�Vc�AE�|�U�G�`hj�"OV���ʎYHib`DU�t�N=�"O  �SO[������ �-y��|(�"O��0���;�m�``�x�~%��"O�$P���GF���ϖ6<@�\��"O�<���sevA�����
��I��y2o��GYF��Ċ��Bq���y�e[=�fِ*�-\�ڨ���ֺ�yrn�Yݾ����@3f�A�,�y⋃�T,%����@D�����	��y�J��@ȸ4�AHȂD���÷b�/�y҇%"���s�E M�l�5F�y����PY6����?CD�5���3�y��Ľ\2<���� "5���;E����y2k��WsD�#��ͣ0i�	Ѕ�8�y��).~���h�	}�\$����y�f�*�j�	W��q���!�ԟ�y�I�[�ZhH��p������Q�y����=�Bd�	o�p�#�ǎ�yBϒMK�򍛸1�8ۢ����y�.V9��ū����rƚ�yRE� :w��j
2m�h�c[��ybA�9Y�n�x߸ޝ��N�-�y� _@�	S�,H�Q�����=�yҊ�g:R� ��8Ek�Uj��y�Ͱ){�p5O't1ƭ�s���y�.��g� �P��1�h��$�y2�#H�V�Ȥ���T���#�y��I5��q��ĄH��]��y�OG�O@���o�w�A���yr
��I?��Ċ�vP�؁��%�y��B�E�����q�Na�q.׳�y`�$&��r`��:�:0��D̊�yr%��;�TP��ӗI ١Q�ނ�y2��	 $| ��%�?&p�!A�O��y�cO�[?`8���T�*SK��y"l�*�|A(�"Y�x�l�P�$��y҆mINd�S��>x)"S!��yr.��Ɓ2bn�)iM>M@�oſ�y�Ȋ�5���1Nѫ6ƪ������y�^L)�%�@�X��R�H�+�y����/4��p�X�M����dj��yBA��� l>	�y�e����y�ƙO3�x��l��1吅3U�<�ym�r����wA�%���ԭ�0�y�AP�2��6!�($��������yr$�F�T2���%��a`���y�̉�J�D;_e�9�	�`�B�	�hN�&M\<O�����H�aC�Ʉ%���u�SRy�yIqgH�(�B�!eBLA�ϊ�fVmc(�"]�\B䉷R��q�������,�*z"B�I�@�6��'�I2���<V"B�I(S=�h�vH�>_��RVaҽ��C䉤q�l8eO|����2L�?��C�	$*��@�ŊWL��k��$�C�ɖHi���5M�/�ހ@E���@�vC�Ȳ��2D�	�͸�˲=-C�	*�&1gi�,�<QA��
�ܡ�� ��� �+2r��XG�NO�̙��"O�t�O�%����ǖ#@�j�#'"OziPf#ȗKp��e&��^�\��0"O�b���#w�>ݸ外!B�L�s"O����\�k �z��/�$��"O���%�xp|���/ۜ4iޕ	�"O��A�ӎK"d��%؛Z�`q6"OVH`%�d��Pcd��xX6H9A"O�YĄ� ���
BOd�e"O�IPdn���@�B��q5�Y�"O��J�/�u�(p���Av �"O8`�w���Zf��(^�%N�a"O��#�Ntk�\q���/�4�c"O��z�JG�k�H��$�\k��h�%"O�����t����dM�2���%"O4�@#�Ȭ-�j��aڿ�,e�F"OZ�c��I;2ɪm鳀-	k�TaU"O�U�����	i�b�OU0hK��"O�U:�/�]��1�lV�%g�-H�"O���R���xg�����Ģ�.�C@"O$|��(C�XqP�=��4�"O�T    �